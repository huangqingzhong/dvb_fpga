--
-- DVB IP
--
-- Copyright 2020 by Suoto <andre820@gmail.com>
--
-- This file is part of the DVB IP.
--
-- DVB IP is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- DVB IP is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with DVB IP.  If not, see <http://www.gnu.org/licenses/>.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.common_pkg.all;

package ldpc_tables_pkg is

  -- From /home/souto/phase4ground/tables/ldpc/dvb/orig/dvb_16200_s2_c10.txt, table is 40x37 (185.0 bytes)
  -- Resource estimation: 3 x 18 kB BRAMs or 2 x 36 kB BRAMs
  type dvb_16200_s2_c10_t is array (39 downto 0) of std_logic_vector(36 downto 0);

  constant DVB_16200_S2_C10_COLUMN_WIDTHS : integer_array_t := (0 => 2, 1 => 2, 2 => 11, 3 => 11, 4 => 11);

  constant DVB_16200_S2_C10 : dvb_16200_s2_c10_t := (
    0 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(0, 2) & to_unsigned(1558, 11) & to_unsigned(712, 11) & to_unsigned(805, 11)),
    1 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(1, 2) & to_unsigned(1450, 11) & to_unsigned(873, 11) & to_unsigned(1337, 11)),
    2 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(2, 2) & to_unsigned(1741, 11) & to_unsigned(1129, 11) & to_unsigned(1184, 11)),
    3 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(3, 2) & to_unsigned(294, 11) & to_unsigned(806, 11) & to_unsigned(1566, 11)),
    4 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(4, 2) & to_unsigned(482, 11) & to_unsigned(605, 11) & to_unsigned(923, 11)),
    5 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 2) & to_unsigned(926, 11) & to_unsigned(1578, 11) & (10 downto 0 => 'U')),
    6 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 2) & to_unsigned(777, 11) & to_unsigned(1374, 11) & (10 downto 0 => 'U')),
    7 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 2) & to_unsigned(608, 11) & to_unsigned(151, 11) & (10 downto 0 => 'U')),
    8 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 2) & to_unsigned(1195, 11) & to_unsigned(210, 11) & (10 downto 0 => 'U')),
    9 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 2) & to_unsigned(1484, 11) & to_unsigned(692, 11) & (10 downto 0 => 'U')),
    10 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 2) & to_unsigned(427, 11) & to_unsigned(488, 11) & (10 downto 0 => 'U')),
    11 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 2) & to_unsigned(828, 11) & to_unsigned(1124, 11) & (10 downto 0 => 'U')),
    12 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 2) & to_unsigned(874, 11) & to_unsigned(1366, 11) & (10 downto 0 => 'U')),
    13 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 2) & to_unsigned(1500, 11) & to_unsigned(835, 11) & (10 downto 0 => 'U')),
    14 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 2) & to_unsigned(1496, 11) & to_unsigned(502, 11) & (10 downto 0 => 'U')),
    15 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 2) & to_unsigned(1006, 11) & to_unsigned(1701, 11) & (10 downto 0 => 'U')),
    16 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 2) & to_unsigned(1155, 11) & to_unsigned(97, 11) & (10 downto 0 => 'U')),
    17 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 2) & to_unsigned(657, 11) & to_unsigned(1403, 11) & (10 downto 0 => 'U')),
    18 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 2) & to_unsigned(1453, 11) & to_unsigned(624, 11) & (10 downto 0 => 'U')),
    19 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 2) & to_unsigned(429, 11) & to_unsigned(1495, 11) & (10 downto 0 => 'U')),
    20 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 2) & to_unsigned(809, 11) & to_unsigned(385, 11) & (10 downto 0 => 'U')),
    21 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 2) & to_unsigned(367, 11) & to_unsigned(151, 11) & (10 downto 0 => 'U')),
    22 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 2) & to_unsigned(1323, 11) & to_unsigned(202, 11) & (10 downto 0 => 'U')),
    23 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 2) & to_unsigned(960, 11) & to_unsigned(318, 11) & (10 downto 0 => 'U')),
    24 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 2) & to_unsigned(1451, 11) & to_unsigned(1039, 11) & (10 downto 0 => 'U')),
    25 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 2) & to_unsigned(1098, 11) & to_unsigned(1722, 11) & (10 downto 0 => 'U')),
    26 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 2) & to_unsigned(1015, 11) & to_unsigned(1428, 11) & (10 downto 0 => 'U')),
    27 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 2) & to_unsigned(1261, 11) & to_unsigned(1564, 11) & (10 downto 0 => 'U')),
    28 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 2) & to_unsigned(544, 11) & to_unsigned(1190, 11) & (10 downto 0 => 'U')),
    29 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 2) & to_unsigned(1472, 11) & to_unsigned(1246, 11) & (10 downto 0 => 'U')),
    30 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 2) & to_unsigned(508, 11) & to_unsigned(630, 11) & (10 downto 0 => 'U')),
    31 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 2) & to_unsigned(421, 11) & to_unsigned(1704, 11) & (10 downto 0 => 'U')),
    32 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 2) & to_unsigned(284, 11) & to_unsigned(898, 11) & (10 downto 0 => 'U')),
    33 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 2) & to_unsigned(392, 11) & to_unsigned(577, 11) & (10 downto 0 => 'U')),
    34 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 2) & to_unsigned(1155, 11) & to_unsigned(556, 11) & (10 downto 0 => 'U')),
    35 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 2) & to_unsigned(631, 11) & to_unsigned(1000, 11) & (10 downto 0 => 'U')),
    36 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 2) & to_unsigned(732, 11) & to_unsigned(1368, 11) & (10 downto 0 => 'U')),
    37 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 2) & to_unsigned(1328, 11) & to_unsigned(329, 11) & (10 downto 0 => 'U')),
    38 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 2) & to_unsigned(1515, 11) & to_unsigned(506, 11) & (10 downto 0 => 'U')),
    39 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 2) & to_unsigned(1104, 11) & to_unsigned(1172, 11) & (10 downto 0 => 'U'))
  );

  -- From /home/souto/phase4ground/tables/ldpc/dvb/orig/dvb_16200_s2_c1_t2_b1.txt, table is 9x171 (192.375 bytes)
  -- Resource estimation: 10 x 18 kB BRAMs or 5 x 36 kB BRAMs
  type dvb_16200_s2_c1_t2_b1_t is array (8 downto 0) of std_logic_vector(170 downto 0);

  constant DVB_16200_S2_C1_T2_B1_COLUMN_WIDTHS : integer_array_t := (0 => 4, 1 => 14, 2 => 14, 3 => 14, 4 => 14, 5 => 13, 6 => 14, 7 => 14, 8 => 14, 9 => 14, 10 => 14, 11 => 14, 12 => 14);

  constant DVB_16200_S2_C1_T2_B1 : dvb_16200_s2_c1_t2_b1_t := (
    0 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(6295, 14) & to_unsigned(9626, 14) & to_unsigned(304, 14) & to_unsigned(7695, 14) & to_unsigned(4839, 13) & to_unsigned(4936, 14) & to_unsigned(1660, 14) & to_unsigned(144, 14) & to_unsigned(11203, 14) & to_unsigned(5567, 14) & to_unsigned(6347, 14) & to_unsigned(12557, 14)),
    1 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(10691, 14) & to_unsigned(4988, 14) & to_unsigned(3859, 14) & to_unsigned(3734, 14) & to_unsigned(3071, 13) & to_unsigned(3494, 14) & to_unsigned(7687, 14) & to_unsigned(10313, 14) & to_unsigned(5964, 14) & to_unsigned(8069, 14) & to_unsigned(8296, 14) & to_unsigned(11090, 14)),
    2 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(10774, 14) & to_unsigned(3613, 14) & to_unsigned(5208, 14) & to_unsigned(11177, 14) & to_unsigned(7676, 13) & to_unsigned(3549, 14) & to_unsigned(8746, 14) & to_unsigned(6583, 14) & to_unsigned(7239, 14) & to_unsigned(12265, 14) & to_unsigned(2674, 14) & to_unsigned(4292, 14)),
    3 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(11869, 14) & to_unsigned(3708, 14) & to_unsigned(5981, 14) & to_unsigned(8718, 14) & to_unsigned(4908, 13) & to_unsigned(10650, 14) & to_unsigned(6805, 14) & to_unsigned(3334, 14) & to_unsigned(2627, 14) & to_unsigned(10461, 14) & to_unsigned(9285, 14) & to_unsigned(11120, 14)),
    4 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7844, 14) & to_unsigned(3079, 14) & to_unsigned(10773, 14) & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    5 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3385, 14) & to_unsigned(10854, 14) & to_unsigned(5747, 14) & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    6 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1360, 14) & to_unsigned(12010, 14) & to_unsigned(12202, 14) & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    7 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6189, 14) & to_unsigned(4241, 14) & to_unsigned(2343, 14) & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    8 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9840, 14) & to_unsigned(12726, 14) & to_unsigned(4977, 14) & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U'))
  );

  -- From /home/souto/phase4ground/tables/ldpc/dvb/orig/dvb_16200_s2_c2_t2_b8.txt, table is 15x170 (318.75 bytes)
  -- Resource estimation: 10 x 18 kB BRAMs or 5 x 36 kB BRAMs
  type dvb_16200_s2_c2_t2_b8_t is array (14 downto 0) of std_logic_vector(169 downto 0);

  constant DVB_16200_S2_C2_T2_B8_COLUMN_WIDTHS : integer_array_t := (0 => 4, 1 => 14, 2 => 14, 3 => 14, 4 => 14, 5 => 14, 6 => 14, 7 => 14, 8 => 13, 9 => 14, 10 => 14, 11 => 14, 12 => 13);

  constant DVB_16200_S2_C2_T2_B8 : dvb_16200_s2_c2_t2_b8_t := (
    0 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(416, 14) & to_unsigned(8909, 14) & to_unsigned(4156, 14) & to_unsigned(3216, 14) & to_unsigned(3112, 14) & to_unsigned(2560, 14) & to_unsigned(2912, 14) & to_unsigned(6405, 13) & to_unsigned(8593, 14) & to_unsigned(4969, 14) & to_unsigned(6723, 14) & to_unsigned(6912, 13)),
    1 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(8978, 14) & to_unsigned(3011, 14) & to_unsigned(4339, 14) & to_unsigned(9312, 14) & to_unsigned(6396, 14) & to_unsigned(2957, 14) & to_unsigned(7288, 14) & to_unsigned(5485, 13) & to_unsigned(6031, 14) & to_unsigned(10218, 14) & to_unsigned(2226, 14) & to_unsigned(3575, 13)),
    2 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(3383, 14) & to_unsigned(10059, 14) & to_unsigned(1114, 14) & to_unsigned(10008, 14) & to_unsigned(10147, 14) & to_unsigned(9384, 14) & to_unsigned(4290, 14) & to_unsigned(434, 13) & to_unsigned(5139, 14) & to_unsigned(3536, 14) & to_unsigned(1965, 14) & to_unsigned(2291, 13)),
    3 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(2797, 14) & to_unsigned(3693, 14) & to_unsigned(7615, 14) & to_unsigned(7077, 14) & to_unsigned(743, 14) & to_unsigned(1941, 14) & to_unsigned(8716, 14) & to_unsigned(6215, 13) & to_unsigned(3840, 14) & to_unsigned(5140, 14) & to_unsigned(4582, 14) & to_unsigned(5420, 13)),
    4 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(6110, 14) & to_unsigned(8551, 14) & to_unsigned(1515, 14) & to_unsigned(7404, 14) & to_unsigned(4879, 14) & to_unsigned(4946, 14) & to_unsigned(5383, 14) & to_unsigned(1831, 13) & to_unsigned(3441, 14) & to_unsigned(9569, 14) & to_unsigned(10472, 14) & to_unsigned(4306, 13)),
    5 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1505, 14) & to_unsigned(5682, 14) & to_unsigned(7778, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U')),
    6 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7172, 14) & to_unsigned(6830, 14) & to_unsigned(6623, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U')),
    7 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7281, 14) & to_unsigned(3941, 14) & to_unsigned(3505, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U')),
    8 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10270, 14) & to_unsigned(8669, 14) & to_unsigned(914, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U')),
    9 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3622, 14) & to_unsigned(7563, 14) & to_unsigned(9388, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U')),
    10 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9930, 14) & to_unsigned(5058, 14) & to_unsigned(4554, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U')),
    11 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4844, 14) & to_unsigned(9609, 14) & to_unsigned(2707, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U')),
    12 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6883, 14) & to_unsigned(3237, 14) & to_unsigned(1714, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U')),
    13 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4768, 14) & to_unsigned(3878, 14) & to_unsigned(10017, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U')),
    14 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10127, 14) & to_unsigned(3334, 14) & to_unsigned(8267, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U'))
  );

  -- From /home/souto/phase4ground/tables/ldpc/dvb/orig/dvb_16200_s2_c3_t2_b9.txt, table is 18x168 (378.0 bytes)
  -- Resource estimation: 10 x 18 kB BRAMs or 5 x 36 kB BRAMs
  type dvb_16200_s2_c3_t2_b9_t is array (17 downto 0) of std_logic_vector(167 downto 0);

  constant DVB_16200_S2_C3_T2_B9_COLUMN_WIDTHS : integer_array_t := (0 => 4, 1 => 14, 2 => 14, 3 => 14, 4 => 14, 5 => 14, 6 => 14, 7 => 13, 8 => 13, 9 => 13, 10 => 14, 11 => 13, 12 => 14);

  constant DVB_16200_S2_C3_T2_B9 : dvb_16200_s2_c3_t2_b9_t := (
    0 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(5650, 14) & to_unsigned(4143, 14) & to_unsigned(8750, 14) & to_unsigned(583, 14) & to_unsigned(6720, 14) & to_unsigned(8071, 14) & to_unsigned(635, 13) & to_unsigned(1767, 13) & to_unsigned(1344, 13) & to_unsigned(6922, 14) & to_unsigned(738, 13) & to_unsigned(6658, 14)),
    1 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(5696, 14) & to_unsigned(1685, 14) & to_unsigned(3207, 14) & to_unsigned(415, 14) & to_unsigned(7019, 14) & to_unsigned(5023, 14) & to_unsigned(5608, 13) & to_unsigned(2605, 13) & to_unsigned(857, 13) & to_unsigned(6915, 14) & to_unsigned(1770, 13) & to_unsigned(8016, 14)),
    2 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(3992, 14) & to_unsigned(771, 14) & to_unsigned(2190, 14) & to_unsigned(7258, 14) & to_unsigned(8970, 14) & to_unsigned(7792, 14) & to_unsigned(1802, 13) & to_unsigned(1866, 13) & to_unsigned(6137, 13) & to_unsigned(8841, 14) & to_unsigned(886, 13) & to_unsigned(1931, 14)),
    3 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(4108, 14) & to_unsigned(3781, 14) & to_unsigned(7577, 14) & to_unsigned(6810, 14) & to_unsigned(9322, 14) & to_unsigned(8226, 14) & to_unsigned(5396, 13) & to_unsigned(5867, 13) & to_unsigned(4428, 13) & to_unsigned(8827, 14) & to_unsigned(7766, 13) & to_unsigned(2254, 14)),
    4 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(4247, 14) & to_unsigned(888, 14) & to_unsigned(4367, 14) & to_unsigned(8821, 14) & to_unsigned(9660, 14) & to_unsigned(324, 14) & to_unsigned(5864, 13) & to_unsigned(4774, 13) & to_unsigned(227, 13) & to_unsigned(7889, 14) & to_unsigned(6405, 13) & to_unsigned(8963, 14)),
    5 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(9693, 14) & to_unsigned(500, 14) & to_unsigned(2520, 14) & to_unsigned(2227, 14) & to_unsigned(1811, 14) & to_unsigned(9330, 14) & to_unsigned(1928, 13) & to_unsigned(5140, 13) & to_unsigned(4030, 13) & to_unsigned(4824, 14) & to_unsigned(806, 13) & to_unsigned(3134, 14)),
    6 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1652, 14) & to_unsigned(8171, 14) & to_unsigned(1435, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U')),
    7 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3366, 14) & to_unsigned(6543, 14) & to_unsigned(3745, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U')),
    8 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9286, 14) & to_unsigned(8509, 14) & to_unsigned(4645, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U')),
    9 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7397, 14) & to_unsigned(5790, 14) & to_unsigned(8972, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U')),
    10 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6597, 14) & to_unsigned(4422, 14) & to_unsigned(1799, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U')),
    11 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9276, 14) & to_unsigned(4041, 14) & to_unsigned(3847, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U')),
    12 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(8683, 14) & to_unsigned(7378, 14) & to_unsigned(4946, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U')),
    13 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5348, 14) & to_unsigned(1993, 14) & to_unsigned(9186, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U')),
    14 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6724, 14) & to_unsigned(9015, 14) & to_unsigned(5646, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U')),
    15 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4502, 14) & to_unsigned(4439, 14) & to_unsigned(8474, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U')),
    16 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5107, 14) & to_unsigned(7342, 14) & to_unsigned(9442, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U')),
    17 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1387, 14) & to_unsigned(8910, 14) & to_unsigned(2660, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U') & (12 downto 0 => 'U') & (13 downto 0 => 'U'))
  );

  -- From /home/souto/phase4ground/tables/ldpc/dvb/orig/dvb_16200_s2_c4_t2_b2.txt, table is 20x100 (250.0 bytes)
  -- Resource estimation: 6 x 18 kB BRAMs or 3 x 36 kB BRAMs
  type dvb_16200_s2_c4_t2_b2_t is array (19 downto 0) of std_logic_vector(99 downto 0);

  constant DVB_16200_S2_C4_T2_B2_COLUMN_WIDTHS : integer_array_t := (0 => 3, 1 => 5, 2 => 14, 3 => 13, 4 => 13, 5 => 13, 6 => 13, 7 => 13, 8 => 13);

  constant DVB_16200_S2_C4_T2_B2 : dvb_16200_s2_c4_t2_b2_t := (
    0 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(20, 5) & to_unsigned(712, 14) & to_unsigned(2386, 13) & to_unsigned(6354, 13) & to_unsigned(4061, 13) & to_unsigned(1062, 13) & to_unsigned(5045, 13) & to_unsigned(5158, 13)),
    1 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(21, 5) & to_unsigned(2543, 14) & to_unsigned(5748, 13) & to_unsigned(4822, 13) & to_unsigned(2348, 13) & to_unsigned(3089, 13) & to_unsigned(6328, 13) & to_unsigned(5876, 13)),
    2 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(22, 5) & to_unsigned(926, 14) & to_unsigned(5701, 13) & to_unsigned(269, 13) & to_unsigned(3693, 13) & to_unsigned(2438, 13) & to_unsigned(3190, 13) & to_unsigned(3507, 13)),
    3 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(23, 5) & to_unsigned(2802, 14) & to_unsigned(4520, 13) & to_unsigned(3577, 13) & to_unsigned(5324, 13) & to_unsigned(1091, 13) & to_unsigned(4667, 13) & to_unsigned(4449, 13)),
    4 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(24, 5) & to_unsigned(5140, 14) & to_unsigned(2003, 13) & to_unsigned(1263, 13) & to_unsigned(4742, 13) & to_unsigned(6497, 13) & to_unsigned(1185, 13) & to_unsigned(6202, 13)),
    5 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(0, 5) & to_unsigned(4046, 14) & to_unsigned(6934, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    6 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(1, 5) & to_unsigned(2855, 14) & to_unsigned(66, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    7 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(2, 5) & to_unsigned(6694, 14) & to_unsigned(212, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    8 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(3, 5) & to_unsigned(3439, 14) & to_unsigned(1158, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    9 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(4, 5) & to_unsigned(3850, 14) & to_unsigned(4422, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    10 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(5, 5) & to_unsigned(5924, 14) & to_unsigned(290, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    11 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(6, 5) & to_unsigned(1467, 14) & to_unsigned(4049, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    12 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(7, 5) & to_unsigned(7820, 14) & to_unsigned(2242, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    13 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(8, 5) & to_unsigned(4606, 14) & to_unsigned(3080, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    14 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(9, 5) & to_unsigned(4633, 14) & to_unsigned(7877, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    15 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(10, 5) & to_unsigned(3884, 14) & to_unsigned(6868, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    16 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(11, 5) & to_unsigned(8935, 14) & to_unsigned(4996, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    17 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(12, 5) & to_unsigned(3028, 14) & to_unsigned(764, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    18 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(13, 5) & to_unsigned(5988, 14) & to_unsigned(1057, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    19 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(14, 5) & to_unsigned(7411, 14) & to_unsigned(3450, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U'))
  );

  -- From /home/souto/phase4ground/tables/ldpc/dvb/orig/dvb_16200_s2_c5.txt, table is 27x160 (540.0 bytes)
  -- Resource estimation: 9 x 18 kB BRAMs or 5 x 36 kB BRAMs
  type dvb_16200_s2_c5_t is array (26 downto 0) of std_logic_vector(159 downto 0);

  constant DVB_16200_S2_C5_COLUMN_WIDTHS : integer_array_t := (0 => 4, 1 => 13, 2 => 13, 3 => 13, 4 => 13, 5 => 13, 6 => 13, 7 => 13, 8 => 13, 9 => 13, 10 => 13, 11 => 13, 12 => 13);

  constant DVB_16200_S2_C5 : dvb_16200_s2_c5_t := (
    0 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(2765, 13) & to_unsigned(5713, 13) & to_unsigned(6426, 13) & to_unsigned(3596, 13) & to_unsigned(1374, 13) & to_unsigned(4811, 13) & to_unsigned(2182, 13) & to_unsigned(544, 13) & to_unsigned(3394, 13) & to_unsigned(2840, 13) & to_unsigned(4310, 13) & to_unsigned(771, 13)),
    1 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(4951, 13) & to_unsigned(211, 13) & to_unsigned(2208, 13) & to_unsigned(723, 13) & to_unsigned(1246, 13) & to_unsigned(2928, 13) & to_unsigned(398, 13) & to_unsigned(5739, 13) & to_unsigned(265, 13) & to_unsigned(5601, 13) & to_unsigned(5993, 13) & to_unsigned(2615, 13)),
    2 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(210, 13) & to_unsigned(4730, 13) & to_unsigned(5777, 13) & to_unsigned(3096, 13) & to_unsigned(4282, 13) & to_unsigned(6238, 13) & to_unsigned(4939, 13) & to_unsigned(1119, 13) & to_unsigned(6463, 13) & to_unsigned(5298, 13) & to_unsigned(6320, 13) & to_unsigned(4016, 13)),
    3 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(4167, 13) & to_unsigned(2063, 13) & to_unsigned(4757, 13) & to_unsigned(3157, 13) & to_unsigned(5664, 13) & to_unsigned(3956, 13) & to_unsigned(6045, 13) & to_unsigned(563, 13) & to_unsigned(4284, 13) & to_unsigned(2441, 13) & to_unsigned(3412, 13) & to_unsigned(6334, 13)),
    4 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(4201, 13) & to_unsigned(2428, 13) & to_unsigned(4474, 13) & to_unsigned(59, 13) & to_unsigned(1721, 13) & to_unsigned(736, 13) & to_unsigned(2997, 13) & to_unsigned(428, 13) & to_unsigned(3807, 13) & to_unsigned(1513, 13) & to_unsigned(4732, 13) & to_unsigned(6195, 13)),
    5 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(2670, 13) & to_unsigned(3081, 13) & to_unsigned(5139, 13) & to_unsigned(3736, 13) & to_unsigned(1999, 13) & to_unsigned(5889, 13) & to_unsigned(4362, 13) & to_unsigned(3806, 13) & to_unsigned(4534, 13) & to_unsigned(5409, 13) & to_unsigned(6384, 13) & to_unsigned(5809, 13)),
    6 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(5516, 13) & to_unsigned(1622, 13) & to_unsigned(2906, 13) & to_unsigned(3285, 13) & to_unsigned(1257, 13) & to_unsigned(5797, 13) & to_unsigned(3816, 13) & to_unsigned(817, 13) & to_unsigned(875, 13) & to_unsigned(2311, 13) & to_unsigned(3543, 13) & to_unsigned(1205, 13)),
    7 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(4244, 13) & to_unsigned(2184, 13) & to_unsigned(5415, 13) & to_unsigned(1705, 13) & to_unsigned(5642, 13) & to_unsigned(4886, 13) & to_unsigned(2333, 13) & to_unsigned(287, 13) & to_unsigned(1848, 13) & to_unsigned(1121, 13) & to_unsigned(3595, 13) & to_unsigned(6022, 13)),
    8 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(2142, 13) & to_unsigned(2830, 13) & to_unsigned(4069, 13) & to_unsigned(5654, 13) & to_unsigned(1295, 13) & to_unsigned(2951, 13) & to_unsigned(3919, 13) & to_unsigned(1356, 13) & to_unsigned(884, 13) & to_unsigned(1786, 13) & to_unsigned(396, 13) & to_unsigned(4738, 13)),
    9 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(0, 13) & to_unsigned(2161, 13) & to_unsigned(2653, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    10 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1, 13) & to_unsigned(1380, 13) & to_unsigned(1461, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    11 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(2, 13) & to_unsigned(2502, 13) & to_unsigned(3707, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    12 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3, 13) & to_unsigned(3971, 13) & to_unsigned(1057, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    13 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 13) & to_unsigned(5985, 13) & to_unsigned(6062, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    14 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 13) & to_unsigned(1733, 13) & to_unsigned(6028, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    15 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 13) & to_unsigned(3786, 13) & to_unsigned(1936, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    16 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 13) & to_unsigned(4292, 13) & to_unsigned(956, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    17 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(8, 13) & to_unsigned(5692, 13) & to_unsigned(3417, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    18 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9, 13) & to_unsigned(266, 13) & to_unsigned(4878, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    19 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10, 13) & to_unsigned(4913, 13) & to_unsigned(3247, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    20 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(11, 13) & to_unsigned(4763, 13) & to_unsigned(3937, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    21 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(12, 13) & to_unsigned(3590, 13) & to_unsigned(2903, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    22 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(13, 13) & to_unsigned(2566, 13) & to_unsigned(4215, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    23 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(14, 13) & to_unsigned(5208, 13) & to_unsigned(4707, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    24 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(15, 13) & to_unsigned(3940, 13) & to_unsigned(3388, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    25 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(16, 13) & to_unsigned(5109, 13) & to_unsigned(4556, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U')),
    26 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(17, 13) & to_unsigned(4908, 13) & to_unsigned(4177, 13) & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U') & (12 downto 0 => 'U'))
  );

  -- From /home/souto/phase4ground/tables/ldpc/dvb/orig/dvb_16200_s2_c6_t2_b4.txt, table is 30x156 (585.0 bytes)
  -- Resource estimation: 9 x 18 kB BRAMs or 5 x 36 kB BRAMs
  type dvb_16200_s2_c6_t2_b4_t is array (29 downto 0) of std_logic_vector(155 downto 0);

  constant DVB_16200_S2_C6_T2_B4_COLUMN_WIDTHS : integer_array_t := (0 => 4, 1 => 4, 2 => 13, 3 => 13, 4 => 12, 5 => 12, 6 => 11, 7 => 12, 8 => 13, 9 => 12, 10 => 13, 11 => 12, 12 => 13, 13 => 12);

  constant DVB_16200_S2_C6_T2_B4 : dvb_16200_s2_c6_t2_b4_t := (
    0 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(0, 4) & to_unsigned(2084, 13) & to_unsigned(1613, 13) & to_unsigned(1548, 12) & to_unsigned(1286, 12) & to_unsigned(1460, 11) & to_unsigned(3196, 12) & to_unsigned(4297, 13) & to_unsigned(2481, 12) & to_unsigned(3369, 13) & to_unsigned(3451, 12) & to_unsigned(4620, 13) & to_unsigned(2622, 12)),
    1 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(1, 4) & to_unsigned(122, 13) & to_unsigned(1516, 13) & to_unsigned(3448, 12) & to_unsigned(2880, 12) & to_unsigned(1407, 11) & to_unsigned(1847, 12) & to_unsigned(3799, 13) & to_unsigned(3529, 12) & to_unsigned(373, 13) & to_unsigned(971, 12) & to_unsigned(4358, 13) & to_unsigned(3108, 12)),
    2 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(2, 4) & to_unsigned(259, 13) & to_unsigned(3399, 13) & to_unsigned(929, 12) & to_unsigned(2650, 12) & to_unsigned(864, 11) & to_unsigned(3996, 12) & to_unsigned(3833, 13) & to_unsigned(107, 12) & to_unsigned(5287, 13) & to_unsigned(164, 12) & to_unsigned(3125, 13) & to_unsigned(2350, 12)),
    3 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3, 4) & to_unsigned(342, 13) & to_unsigned(3529, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    4 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 4) & to_unsigned(4198, 13) & to_unsigned(2147, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    5 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 4) & to_unsigned(1880, 13) & to_unsigned(4836, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    6 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 4) & to_unsigned(3864, 13) & to_unsigned(4910, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    7 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 4) & to_unsigned(243, 13) & to_unsigned(1542, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    8 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(8, 4) & to_unsigned(3011, 13) & to_unsigned(1436, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    9 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9, 4) & to_unsigned(2167, 13) & to_unsigned(2512, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    10 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10, 4) & to_unsigned(4606, 13) & to_unsigned(1003, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    11 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(11, 4) & to_unsigned(2835, 13) & to_unsigned(705, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    12 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(12, 4) & to_unsigned(3426, 13) & to_unsigned(2365, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    13 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(13, 4) & to_unsigned(3848, 13) & to_unsigned(2474, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    14 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(14, 4) & to_unsigned(1360, 13) & to_unsigned(1743, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    15 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(0, 4) & to_unsigned(163, 13) & to_unsigned(2536, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    16 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1, 4) & to_unsigned(2583, 13) & to_unsigned(1180, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    17 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(2, 4) & to_unsigned(1542, 13) & to_unsigned(509, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    18 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3, 4) & to_unsigned(4418, 13) & to_unsigned(1005, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    19 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 4) & to_unsigned(5212, 13) & to_unsigned(5117, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    20 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 4) & to_unsigned(2155, 13) & to_unsigned(2922, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    21 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 4) & to_unsigned(347, 13) & to_unsigned(2696, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    22 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 4) & to_unsigned(226, 13) & to_unsigned(4296, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    23 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(8, 4) & to_unsigned(1560, 13) & to_unsigned(487, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    24 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9, 4) & to_unsigned(3926, 13) & to_unsigned(1640, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    25 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10, 4) & to_unsigned(149, 13) & to_unsigned(2928, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    26 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(11, 4) & to_unsigned(2364, 13) & to_unsigned(563, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    27 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(12, 4) & to_unsigned(635, 13) & to_unsigned(688, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    28 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(13, 4) & to_unsigned(231, 13) & to_unsigned(1684, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U')),
    29 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(14, 4) & to_unsigned(1129, 13) & to_unsigned(3894, 13) & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U') & (12 downto 0 => 'U') & (11 downto 0 => 'U'))
  );

  -- From /home/souto/phase4ground/tables/ldpc/dvb/orig/dvb_16200_s2_c7_t2_b5.txt, table is 33x133 (548.625 bytes)
  -- Resource estimation: 8 x 18 kB BRAMs or 4 x 36 kB BRAMs
  type dvb_16200_s2_c7_t2_b5_t is array (32 downto 0) of std_logic_vector(132 downto 0);

  constant DVB_16200_S2_C7_T2_B5_COLUMN_WIDTHS : integer_array_t := (0 => 4, 1 => 4, 2 => 13, 3 => 12, 4 => 13, 5 => 11, 6 => 10, 7 => 12, 8 => 11, 9 => 12, 10 => 10, 11 => 10, 12 => 11);

  constant DVB_16200_S2_C7_T2_B5 : dvb_16200_s2_c7_t2_b5_t := (
    0 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(3, 4) & to_unsigned(3198, 13) & to_unsigned(478, 12) & to_unsigned(4207, 13) & to_unsigned(1481, 11) & to_unsigned(1009, 10) & to_unsigned(2616, 12) & to_unsigned(1924, 11) & to_unsigned(3437, 12) & to_unsigned(554, 10) & to_unsigned(683, 10) & to_unsigned(1801, 11)),
    1 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 4) & to_unsigned(2681, 13) & to_unsigned(2135, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    2 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 4) & to_unsigned(3107, 13) & to_unsigned(4027, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    3 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 4) & to_unsigned(2637, 13) & to_unsigned(3373, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    4 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 4) & to_unsigned(3830, 13) & to_unsigned(3449, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    5 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(8, 4) & to_unsigned(4129, 13) & to_unsigned(2060, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    6 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9, 4) & to_unsigned(4184, 13) & to_unsigned(2742, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    7 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10, 4) & to_unsigned(3946, 13) & to_unsigned(1070, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    8 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(11, 4) & to_unsigned(2239, 13) & to_unsigned(984, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    9 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(0, 4) & to_unsigned(1458, 13) & to_unsigned(3031, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    10 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1, 4) & to_unsigned(3003, 13) & to_unsigned(1328, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    11 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(2, 4) & to_unsigned(1137, 13) & to_unsigned(1716, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    12 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3, 4) & to_unsigned(132, 13) & to_unsigned(3725, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    13 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 4) & to_unsigned(1817, 13) & to_unsigned(638, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    14 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 4) & to_unsigned(1774, 13) & to_unsigned(3447, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    15 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 4) & to_unsigned(3632, 13) & to_unsigned(1257, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    16 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 4) & to_unsigned(542, 13) & to_unsigned(3694, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    17 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(8, 4) & to_unsigned(1015, 13) & to_unsigned(1945, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    18 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9, 4) & to_unsigned(1948, 13) & to_unsigned(412, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    19 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10, 4) & to_unsigned(995, 13) & to_unsigned(2238, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    20 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(11, 4) & to_unsigned(4141, 13) & to_unsigned(1907, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    21 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(0, 4) & to_unsigned(2480, 13) & to_unsigned(3079, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    22 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1, 4) & to_unsigned(3021, 13) & to_unsigned(1088, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    23 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(2, 4) & to_unsigned(713, 13) & to_unsigned(1379, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    24 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3, 4) & to_unsigned(997, 13) & to_unsigned(3903, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    25 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 4) & to_unsigned(2323, 13) & to_unsigned(3361, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    26 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 4) & to_unsigned(1110, 13) & to_unsigned(986, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    27 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 4) & to_unsigned(2532, 13) & to_unsigned(142, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    28 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 4) & to_unsigned(1690, 13) & to_unsigned(2405, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    29 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(8, 4) & to_unsigned(1298, 13) & to_unsigned(1881, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    30 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9, 4) & to_unsigned(615, 13) & to_unsigned(174, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    31 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10, 4) & to_unsigned(1648, 13) & to_unsigned(3112, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U')),
    32 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(11, 4) & to_unsigned(1415, 13) & to_unsigned(2808, 12) & (12 downto 0 => 'U') & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U'))
  );

  -- From /home/souto/phase4ground/tables/ldpc/dvb/orig/dvb_16200_s2_c8_t2_b6.txt, table is 35x30 (131.25 bytes)
  -- Resource estimation: 2 x 18 kB BRAMs or 1 x 36 kB BRAMs
  type dvb_16200_s2_c8_t2_b6_t is array (34 downto 0) of std_logic_vector(29 downto 0);

  constant DVB_16200_S2_C8_T2_B6_COLUMN_WIDTHS : integer_array_t := (0 => 2, 1 => 4, 2 => 12, 3 => 12);

  constant DVB_16200_S2_C8_T2_B6 : dvb_16200_s2_c8_t2_b6_t := (
    0 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(5, 4) & to_unsigned(896, 12) & to_unsigned(1565, 12)),
    1 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(6, 4) & to_unsigned(2493, 12) & to_unsigned(184, 12)),
    2 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(7, 4) & to_unsigned(212, 12) & to_unsigned(3210, 12)),
    3 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(8, 4) & to_unsigned(727, 12) & to_unsigned(1339, 12)),
    4 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(9, 4) & to_unsigned(3428, 12) & to_unsigned(612, 12)),
    5 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 4) & to_unsigned(2663, 12) & to_unsigned(1947, 12)),
    6 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 4) & to_unsigned(230, 12) & to_unsigned(2695, 12)),
    7 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 4) & to_unsigned(2025, 12) & to_unsigned(2794, 12)),
    8 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 4) & to_unsigned(3039, 12) & to_unsigned(283, 12)),
    9 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 4) & to_unsigned(862, 12) & to_unsigned(2889, 12)),
    10 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(5, 4) & to_unsigned(376, 12) & to_unsigned(2110, 12)),
    11 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(6, 4) & to_unsigned(2034, 12) & to_unsigned(2286, 12)),
    12 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(7, 4) & to_unsigned(951, 12) & to_unsigned(2068, 12)),
    13 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(8, 4) & to_unsigned(3108, 12) & to_unsigned(3542, 12)),
    14 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(9, 4) & to_unsigned(307, 12) & to_unsigned(1421, 12)),
    15 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 4) & to_unsigned(2272, 12) & to_unsigned(1197, 12)),
    16 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 4) & to_unsigned(1800, 12) & to_unsigned(3280, 12)),
    17 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 4) & to_unsigned(331, 12) & to_unsigned(2308, 12)),
    18 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 4) & to_unsigned(465, 12) & to_unsigned(2552, 12)),
    19 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 4) & to_unsigned(1038, 12) & to_unsigned(2479, 12)),
    20 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(5, 4) & to_unsigned(1383, 12) & to_unsigned(343, 12)),
    21 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(6, 4) & to_unsigned(94, 12) & to_unsigned(236, 12)),
    22 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(7, 4) & to_unsigned(2619, 12) & to_unsigned(121, 12)),
    23 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(8, 4) & to_unsigned(1497, 12) & to_unsigned(2774, 12)),
    24 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(9, 4) & to_unsigned(2116, 12) & to_unsigned(1855, 12)),
    25 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 4) & to_unsigned(722, 12) & to_unsigned(1584, 12)),
    26 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 4) & to_unsigned(2767, 12) & to_unsigned(1881, 12)),
    27 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 4) & to_unsigned(2701, 12) & to_unsigned(1610, 12)),
    28 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 4) & to_unsigned(3283, 12) & to_unsigned(1732, 12)),
    29 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 4) & to_unsigned(168, 12) & to_unsigned(1099, 12)),
    30 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(5, 4) & to_unsigned(3074, 12) & to_unsigned(243, 12)),
    31 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(6, 4) & to_unsigned(3460, 12) & to_unsigned(945, 12)),
    32 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(7, 4) & to_unsigned(2049, 12) & to_unsigned(1746, 12)),
    33 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(8, 4) & to_unsigned(566, 12) & to_unsigned(1427, 12)),
    34 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(9, 4) & to_unsigned(3545, 12) & to_unsigned(1168, 12))
  );

  -- From /home/souto/phase4ground/tables/ldpc/dvb/orig/dvb_16200_s2_c9_t2_b7.txt, table is 37x139 (642.875 bytes)
  -- Resource estimation: 8 x 18 kB BRAMs or 4 x 36 kB BRAMs
  type dvb_16200_s2_c9_t2_b7_t is array (36 downto 0) of std_logic_vector(138 downto 0);

  constant DVB_16200_S2_C9_T2_B7_COLUMN_WIDTHS : integer_array_t := (0 => 4, 1 => 3, 2 => 12, 3 => 12, 4 => 11, 5 => 10, 6 => 10, 7 => 10, 8 => 11, 9 => 9, 10 => 12, 11 => 12, 12 => 11, 13 => 12);

  constant DVB_16200_S2_C9_T2_B7 : dvb_16200_s2_c9_t2_b7_t := (
    0 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(3, 3) & to_unsigned(2409, 12) & to_unsigned(499, 12) & to_unsigned(1481, 11) & to_unsigned(908, 10) & to_unsigned(559, 10) & to_unsigned(716, 10) & to_unsigned(1270, 11) & to_unsigned(333, 9) & to_unsigned(2508, 12) & to_unsigned(2264, 12) & to_unsigned(1702, 11) & to_unsigned(2805, 12)),
    1 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 3) & to_unsigned(2447, 12) & to_unsigned(1926, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    2 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 3) & to_unsigned(414, 12) & to_unsigned(1224, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    3 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 3) & to_unsigned(2114, 12) & to_unsigned(842, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    4 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 3) & to_unsigned(212, 12) & to_unsigned(573, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    5 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(0, 3) & to_unsigned(2383, 12) & to_unsigned(2112, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    6 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1, 3) & to_unsigned(2286, 12) & to_unsigned(2348, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    7 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(2, 3) & to_unsigned(545, 12) & to_unsigned(819, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    8 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3, 3) & to_unsigned(1264, 12) & to_unsigned(143, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    9 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 3) & to_unsigned(1701, 12) & to_unsigned(2258, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    10 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 3) & to_unsigned(964, 12) & to_unsigned(166, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    11 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 3) & to_unsigned(114, 12) & to_unsigned(2413, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    12 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 3) & to_unsigned(2243, 12) & to_unsigned(81, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    13 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(0, 3) & to_unsigned(1245, 12) & to_unsigned(1581, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    14 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1, 3) & to_unsigned(775, 12) & to_unsigned(169, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    15 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(2, 3) & to_unsigned(1696, 12) & to_unsigned(1104, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    16 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3, 3) & to_unsigned(1914, 12) & to_unsigned(2831, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    17 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 3) & to_unsigned(532, 12) & to_unsigned(1450, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    18 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 3) & to_unsigned(91, 12) & to_unsigned(974, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    19 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 3) & to_unsigned(497, 12) & to_unsigned(2228, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    20 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 3) & to_unsigned(2326, 12) & to_unsigned(1579, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    21 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(0, 3) & to_unsigned(2482, 12) & to_unsigned(256, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    22 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1, 3) & to_unsigned(1117, 12) & to_unsigned(1261, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    23 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(2, 3) & to_unsigned(1257, 12) & to_unsigned(1658, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    24 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3, 3) & to_unsigned(1478, 12) & to_unsigned(1225, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    25 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 3) & to_unsigned(2511, 12) & to_unsigned(980, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    26 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 3) & to_unsigned(2320, 12) & to_unsigned(2675, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    27 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 3) & to_unsigned(435, 12) & to_unsigned(1278, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    28 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 3) & to_unsigned(228, 12) & to_unsigned(503, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    29 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(0, 3) & to_unsigned(1885, 12) & to_unsigned(2369, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    30 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1, 3) & to_unsigned(57, 12) & to_unsigned(483, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    31 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(2, 3) & to_unsigned(838, 12) & to_unsigned(1050, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    32 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3, 3) & to_unsigned(1231, 12) & to_unsigned(1990, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    33 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 3) & to_unsigned(1738, 12) & to_unsigned(68, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    34 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 3) & to_unsigned(2392, 12) & to_unsigned(951, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    35 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 3) & to_unsigned(163, 12) & to_unsigned(645, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U')),
    36 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 3) & to_unsigned(2644, 12) & to_unsigned(1704, 12) & (10 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (9 downto 0 => 'U') & (10 downto 0 => 'U') & (8 downto 0 => 'U') & (11 downto 0 => 'U') & (11 downto 0 => 'U') & (10 downto 0 => 'U') & (11 downto 0 => 'U'))
  );

  -- From /home/souto/phase4ground/tables/ldpc/dvb/orig/dvb_64800_s2_b1.txt, table is 45x196 (1102.5 bytes)
  -- Resource estimation: 11 x 18 kB BRAMs or 6 x 36 kB BRAMs
  type dvb_64800_s2_b1_t is array (44 downto 0) of std_logic_vector(195 downto 0);

  constant DVB_64800_S2_B1_COLUMN_WIDTHS : integer_array_t := (0 => 4, 1 => 16, 2 => 16, 3 => 16, 4 => 16, 5 => 16, 6 => 16, 7 => 16, 8 => 16, 9 => 16, 10 => 16, 11 => 16, 12 => 16);

  constant DVB_64800_S2_B1 : dvb_64800_s2_b1_t := (
    0 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(23606, 16) & to_unsigned(36098, 16) & to_unsigned(1140, 16) & to_unsigned(28859, 16) & to_unsigned(18148, 16) & to_unsigned(18510, 16) & to_unsigned(6226, 16) & to_unsigned(540, 16) & to_unsigned(42014, 16) & to_unsigned(20879, 16) & to_unsigned(23802, 16) & to_unsigned(47088, 16)),
    1 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(16419, 16) & to_unsigned(24928, 16) & to_unsigned(16609, 16) & to_unsigned(17248, 16) & to_unsigned(7693, 16) & to_unsigned(24997, 16) & to_unsigned(42587, 16) & to_unsigned(16858, 16) & to_unsigned(34921, 16) & to_unsigned(21042, 16) & to_unsigned(37024, 16) & to_unsigned(20692, 16)),
    2 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(1874, 16) & to_unsigned(40094, 16) & to_unsigned(18704, 16) & to_unsigned(14474, 16) & to_unsigned(14004, 16) & to_unsigned(11519, 16) & to_unsigned(13106, 16) & to_unsigned(28826, 16) & to_unsigned(38669, 16) & to_unsigned(22363, 16) & to_unsigned(30255, 16) & to_unsigned(31105, 16)),
    3 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(22254, 16) & to_unsigned(40564, 16) & to_unsigned(22645, 16) & to_unsigned(22532, 16) & to_unsigned(6134, 16) & to_unsigned(9176, 16) & to_unsigned(39998, 16) & to_unsigned(23892, 16) & to_unsigned(8937, 16) & to_unsigned(15608, 16) & to_unsigned(16854, 16) & to_unsigned(31009, 16)),
    4 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(8037, 16) & to_unsigned(40401, 16) & to_unsigned(13550, 16) & to_unsigned(19526, 16) & to_unsigned(41902, 16) & to_unsigned(28782, 16) & to_unsigned(13304, 16) & to_unsigned(32796, 16) & to_unsigned(24679, 16) & to_unsigned(27140, 16) & to_unsigned(45980, 16) & to_unsigned(10021, 16)),
    5 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(40540, 16) & to_unsigned(44498, 16) & to_unsigned(13911, 16) & to_unsigned(22435, 16) & to_unsigned(32701, 16) & to_unsigned(18405, 16) & to_unsigned(39929, 16) & to_unsigned(25521, 16) & to_unsigned(12497, 16) & to_unsigned(9851, 16) & to_unsigned(39223, 16) & to_unsigned(34823, 16)),
    6 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(15233, 16) & to_unsigned(45333, 16) & to_unsigned(5041, 16) & to_unsigned(44979, 16) & to_unsigned(45710, 16) & to_unsigned(42150, 16) & to_unsigned(19416, 16) & to_unsigned(1892, 16) & to_unsigned(23121, 16) & to_unsigned(15860, 16) & to_unsigned(8832, 16) & to_unsigned(10308, 16)),
    7 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(10468, 16) & to_unsigned(44296, 16) & to_unsigned(3611, 16) & to_unsigned(1480, 16) & to_unsigned(37581, 16) & to_unsigned(32254, 16) & to_unsigned(13817, 16) & to_unsigned(6883, 16) & to_unsigned(32892, 16) & to_unsigned(40258, 16) & to_unsigned(46538, 16) & to_unsigned(11940, 16)),
    8 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(6705, 16) & to_unsigned(21634, 16) & to_unsigned(28150, 16) & to_unsigned(43757, 16) & to_unsigned(895, 16) & to_unsigned(6547, 16) & to_unsigned(20970, 16) & to_unsigned(28914, 16) & to_unsigned(30117, 16) & to_unsigned(25736, 16) & to_unsigned(41734, 16) & to_unsigned(11392, 16)),
    9 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(22002, 16) & to_unsigned(5739, 16) & to_unsigned(27210, 16) & to_unsigned(27828, 16) & to_unsigned(34192, 16) & to_unsigned(37992, 16) & to_unsigned(10915, 16) & to_unsigned(6998, 16) & to_unsigned(3824, 16) & to_unsigned(42130, 16) & to_unsigned(4494, 16) & to_unsigned(35739, 16)),
    10 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(8515, 16) & to_unsigned(1191, 16) & to_unsigned(13642, 16) & to_unsigned(30950, 16) & to_unsigned(25943, 16) & to_unsigned(12673, 16) & to_unsigned(16726, 16) & to_unsigned(34261, 16) & to_unsigned(31828, 16) & to_unsigned(3340, 16) & to_unsigned(8747, 16) & to_unsigned(39225, 16)),
    11 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(18979, 16) & to_unsigned(17058, 16) & to_unsigned(43130, 16) & to_unsigned(4246, 16) & to_unsigned(4793, 16) & to_unsigned(44030, 16) & to_unsigned(19454, 16) & to_unsigned(29511, 16) & to_unsigned(47929, 16) & to_unsigned(15174, 16) & to_unsigned(24333, 16) & to_unsigned(19354, 16)),
    12 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(16694, 16) & to_unsigned(8381, 16) & to_unsigned(29642, 16) & to_unsigned(46516, 16) & to_unsigned(32224, 16) & to_unsigned(26344, 16) & to_unsigned(9405, 16) & to_unsigned(18292, 16) & to_unsigned(12437, 16) & to_unsigned(27316, 16) & to_unsigned(35466, 16) & to_unsigned(41992, 16)),
    13 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(15642, 16) & to_unsigned(5871, 16) & to_unsigned(46489, 16) & to_unsigned(26723, 16) & to_unsigned(23396, 16) & to_unsigned(7257, 16) & to_unsigned(8974, 16) & to_unsigned(3156, 16) & to_unsigned(37420, 16) & to_unsigned(44823, 16) & to_unsigned(35423, 16) & to_unsigned(13541, 16)),
    14 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(42858, 16) & to_unsigned(32008, 16) & to_unsigned(41282, 16) & to_unsigned(38773, 16) & to_unsigned(26570, 16) & to_unsigned(2702, 16) & to_unsigned(27260, 16) & to_unsigned(46974, 16) & to_unsigned(1469, 16) & to_unsigned(20887, 16) & to_unsigned(27426, 16) & to_unsigned(38553, 16)),
    15 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(22152, 16) & to_unsigned(24261, 16) & to_unsigned(8297, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    16 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(19347, 16) & to_unsigned(9978, 16) & to_unsigned(27802, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    17 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(34991, 16) & to_unsigned(6354, 16) & to_unsigned(33561, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    18 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(29782, 16) & to_unsigned(30875, 16) & to_unsigned(29523, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    19 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9278, 16) & to_unsigned(48512, 16) & to_unsigned(14349, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    20 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(38061, 16) & to_unsigned(4165, 16) & to_unsigned(43878, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    21 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(8548, 16) & to_unsigned(33172, 16) & to_unsigned(34410, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    22 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(22535, 16) & to_unsigned(28811, 16) & to_unsigned(23950, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    23 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(20439, 16) & to_unsigned(4027, 16) & to_unsigned(24186, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    24 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(38618, 16) & to_unsigned(8187, 16) & to_unsigned(30947, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    25 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(35538, 16) & to_unsigned(43880, 16) & to_unsigned(21459, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    26 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7091, 16) & to_unsigned(45616, 16) & to_unsigned(15063, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    27 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5505, 16) & to_unsigned(9315, 16) & to_unsigned(21908, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    28 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(36046, 16) & to_unsigned(32914, 16) & to_unsigned(11836, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    29 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7304, 16) & to_unsigned(39782, 16) & to_unsigned(33721, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    30 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(16905, 16) & to_unsigned(29962, 16) & to_unsigned(12980, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    31 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(11171, 16) & to_unsigned(23709, 16) & to_unsigned(22460, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    32 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(34541, 16) & to_unsigned(9937, 16) & to_unsigned(44500, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    33 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(14035, 16) & to_unsigned(47316, 16) & to_unsigned(8815, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    34 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(15057, 16) & to_unsigned(45482, 16) & to_unsigned(24461, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    35 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(30518, 16) & to_unsigned(36877, 16) & to_unsigned(879, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    36 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7583, 16) & to_unsigned(13364, 16) & to_unsigned(24332, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    37 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(448, 16) & to_unsigned(27056, 16) & to_unsigned(4682, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    38 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(12083, 16) & to_unsigned(31378, 16) & to_unsigned(21670, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    39 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1159, 16) & to_unsigned(18031, 16) & to_unsigned(2221, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    40 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(17028, 16) & to_unsigned(38715, 16) & to_unsigned(9350, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    41 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(17343, 16) & to_unsigned(24530, 16) & to_unsigned(29574, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    42 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(46128, 16) & to_unsigned(31039, 16) & to_unsigned(32818, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    43 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(20373, 16) & to_unsigned(36967, 16) & to_unsigned(18345, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    44 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(46685, 16) & to_unsigned(20622, 16) & to_unsigned(32806, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U'))
  );

  -- From /home/souto/phase4ground/tables/ldpc/dvb/orig/dvb_64800_s2_b10.txt, table is 160x46 (920.0 bytes)
  -- Resource estimation: 3 x 18 kB BRAMs or 2 x 36 kB BRAMs
  type dvb_64800_s2_b10_t is array (159 downto 0) of std_logic_vector(45 downto 0);

  constant DVB_64800_S2_B10_COLUMN_WIDTHS : integer_array_t := (0 => 2, 1 => 5, 2 => 13, 3 => 13, 4 => 13);

  constant DVB_64800_S2_B10 : dvb_64800_s2_b10_t := (
    0 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(0, 5) & to_unsigned(6235, 13) & to_unsigned(2848, 13) & to_unsigned(3222, 13)),
    1 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(1, 5) & to_unsigned(5800, 13) & to_unsigned(3492, 13) & to_unsigned(5348, 13)),
    2 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(2, 5) & to_unsigned(2757, 13) & to_unsigned(927, 13) & to_unsigned(90, 13)),
    3 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(3, 5) & to_unsigned(6961, 13) & to_unsigned(4516, 13) & to_unsigned(4739, 13)),
    4 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(4, 5) & to_unsigned(1172, 13) & to_unsigned(3237, 13) & to_unsigned(6264, 13)),
    5 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(5, 5) & to_unsigned(1927, 13) & to_unsigned(2425, 13) & to_unsigned(3683, 13)),
    6 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(6, 5) & to_unsigned(3714, 13) & to_unsigned(6309, 13) & to_unsigned(2495, 13)),
    7 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(7, 5) & to_unsigned(3070, 13) & to_unsigned(6342, 13) & to_unsigned(7154, 13)),
    8 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(8, 5) & to_unsigned(2428, 13) & to_unsigned(613, 13) & to_unsigned(3761, 13)),
    9 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(9, 5) & to_unsigned(2906, 13) & to_unsigned(264, 13) & to_unsigned(5927, 13)),
    10 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(10, 5) & to_unsigned(1716, 13) & to_unsigned(1950, 13) & to_unsigned(4273, 13)),
    11 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(11, 5) & to_unsigned(4613, 13) & to_unsigned(6179, 13) & to_unsigned(3491, 13)),
    12 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(12, 5) & to_unsigned(4865, 13) & to_unsigned(3286, 13) & to_unsigned(6005, 13)),
    13 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(13, 5) & to_unsigned(1343, 13) & to_unsigned(5923, 13) & to_unsigned(3529, 13)),
    14 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(14, 5) & to_unsigned(4589, 13) & to_unsigned(4035, 13) & to_unsigned(2132, 13)),
    15 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(15, 5) & to_unsigned(1579, 13) & to_unsigned(3920, 13) & to_unsigned(6737, 13)),
    16 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(16, 5) & to_unsigned(1644, 13) & to_unsigned(1191, 13) & to_unsigned(5998, 13)),
    17 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(17, 5) & to_unsigned(1482, 13) & to_unsigned(2381, 13) & to_unsigned(4620, 13)),
    18 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(18, 5) & to_unsigned(6791, 13) & to_unsigned(6014, 13) & to_unsigned(6596, 13)),
    19 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(19, 5) & to_unsigned(2738, 13) & to_unsigned(5918, 13) & to_unsigned(3786, 13)),
    20 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 5) & to_unsigned(5156, 13) & to_unsigned(6166, 13) & (12 downto 0 => 'U')),
    21 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 5) & to_unsigned(1504, 13) & to_unsigned(4356, 13) & (12 downto 0 => 'U')),
    22 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 5) & to_unsigned(130, 13) & to_unsigned(1904, 13) & (12 downto 0 => 'U')),
    23 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 5) & to_unsigned(6027, 13) & to_unsigned(3187, 13) & (12 downto 0 => 'U')),
    24 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 5) & to_unsigned(6718, 13) & to_unsigned(759, 13) & (12 downto 0 => 'U')),
    25 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(5, 5) & to_unsigned(6240, 13) & to_unsigned(2870, 13) & (12 downto 0 => 'U')),
    26 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(6, 5) & to_unsigned(2343, 13) & to_unsigned(1311, 13) & (12 downto 0 => 'U')),
    27 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(7, 5) & to_unsigned(1039, 13) & to_unsigned(5465, 13) & (12 downto 0 => 'U')),
    28 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(8, 5) & to_unsigned(6617, 13) & to_unsigned(2513, 13) & (12 downto 0 => 'U')),
    29 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(9, 5) & to_unsigned(1588, 13) & to_unsigned(5222, 13) & (12 downto 0 => 'U')),
    30 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(10, 5) & to_unsigned(6561, 13) & to_unsigned(535, 13) & (12 downto 0 => 'U')),
    31 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(11, 5) & to_unsigned(4765, 13) & to_unsigned(2054, 13) & (12 downto 0 => 'U')),
    32 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(12, 5) & to_unsigned(5966, 13) & to_unsigned(6892, 13) & (12 downto 0 => 'U')),
    33 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(13, 5) & to_unsigned(1969, 13) & to_unsigned(3869, 13) & (12 downto 0 => 'U')),
    34 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(14, 5) & to_unsigned(3571, 13) & to_unsigned(2420, 13) & (12 downto 0 => 'U')),
    35 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(15, 5) & to_unsigned(4632, 13) & to_unsigned(981, 13) & (12 downto 0 => 'U')),
    36 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(16, 5) & to_unsigned(3215, 13) & to_unsigned(4163, 13) & (12 downto 0 => 'U')),
    37 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(17, 5) & to_unsigned(973, 13) & to_unsigned(3117, 13) & (12 downto 0 => 'U')),
    38 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(18, 5) & to_unsigned(3802, 13) & to_unsigned(6198, 13) & (12 downto 0 => 'U')),
    39 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(19, 5) & to_unsigned(3794, 13) & to_unsigned(3948, 13) & (12 downto 0 => 'U')),
    40 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 5) & to_unsigned(3196, 13) & to_unsigned(6126, 13) & (12 downto 0 => 'U')),
    41 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 5) & to_unsigned(573, 13) & to_unsigned(1909, 13) & (12 downto 0 => 'U')),
    42 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 5) & to_unsigned(850, 13) & to_unsigned(4034, 13) & (12 downto 0 => 'U')),
    43 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 5) & to_unsigned(5622, 13) & to_unsigned(1601, 13) & (12 downto 0 => 'U')),
    44 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 5) & to_unsigned(6005, 13) & to_unsigned(524, 13) & (12 downto 0 => 'U')),
    45 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(5, 5) & to_unsigned(5251, 13) & to_unsigned(5783, 13) & (12 downto 0 => 'U')),
    46 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(6, 5) & to_unsigned(172, 13) & to_unsigned(2032, 13) & (12 downto 0 => 'U')),
    47 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(7, 5) & to_unsigned(1875, 13) & to_unsigned(2475, 13) & (12 downto 0 => 'U')),
    48 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(8, 5) & to_unsigned(497, 13) & to_unsigned(1291, 13) & (12 downto 0 => 'U')),
    49 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(9, 5) & to_unsigned(2566, 13) & to_unsigned(3430, 13) & (12 downto 0 => 'U')),
    50 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(10, 5) & to_unsigned(1249, 13) & to_unsigned(740, 13) & (12 downto 0 => 'U')),
    51 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(11, 5) & to_unsigned(2944, 13) & to_unsigned(1948, 13) & (12 downto 0 => 'U')),
    52 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(12, 5) & to_unsigned(6528, 13) & to_unsigned(2899, 13) & (12 downto 0 => 'U')),
    53 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(13, 5) & to_unsigned(2243, 13) & to_unsigned(3616, 13) & (12 downto 0 => 'U')),
    54 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(14, 5) & to_unsigned(867, 13) & to_unsigned(3733, 13) & (12 downto 0 => 'U')),
    55 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(15, 5) & to_unsigned(1374, 13) & to_unsigned(4702, 13) & (12 downto 0 => 'U')),
    56 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(16, 5) & to_unsigned(4698, 13) & to_unsigned(2285, 13) & (12 downto 0 => 'U')),
    57 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(17, 5) & to_unsigned(4760, 13) & to_unsigned(3917, 13) & (12 downto 0 => 'U')),
    58 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(18, 5) & to_unsigned(1859, 13) & to_unsigned(4058, 13) & (12 downto 0 => 'U')),
    59 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(19, 5) & to_unsigned(6141, 13) & to_unsigned(3527, 13) & (12 downto 0 => 'U')),
    60 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 5) & to_unsigned(2148, 13) & to_unsigned(5066, 13) & (12 downto 0 => 'U')),
    61 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 5) & to_unsigned(1306, 13) & to_unsigned(145, 13) & (12 downto 0 => 'U')),
    62 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 5) & to_unsigned(2319, 13) & to_unsigned(871, 13) & (12 downto 0 => 'U')),
    63 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 5) & to_unsigned(3463, 13) & to_unsigned(1061, 13) & (12 downto 0 => 'U')),
    64 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 5) & to_unsigned(5554, 13) & to_unsigned(6647, 13) & (12 downto 0 => 'U')),
    65 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(5, 5) & to_unsigned(5837, 13) & to_unsigned(339, 13) & (12 downto 0 => 'U')),
    66 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(6, 5) & to_unsigned(5821, 13) & to_unsigned(4932, 13) & (12 downto 0 => 'U')),
    67 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(7, 5) & to_unsigned(6356, 13) & to_unsigned(4756, 13) & (12 downto 0 => 'U')),
    68 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(8, 5) & to_unsigned(3930, 13) & to_unsigned(418, 13) & (12 downto 0 => 'U')),
    69 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(9, 5) & to_unsigned(211, 13) & to_unsigned(3094, 13) & (12 downto 0 => 'U')),
    70 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(10, 5) & to_unsigned(1007, 13) & to_unsigned(4928, 13) & (12 downto 0 => 'U')),
    71 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(11, 5) & to_unsigned(3584, 13) & to_unsigned(1235, 13) & (12 downto 0 => 'U')),
    72 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(12, 5) & to_unsigned(6982, 13) & to_unsigned(2869, 13) & (12 downto 0 => 'U')),
    73 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(13, 5) & to_unsigned(1612, 13) & to_unsigned(1013, 13) & (12 downto 0 => 'U')),
    74 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(14, 5) & to_unsigned(953, 13) & to_unsigned(4964, 13) & (12 downto 0 => 'U')),
    75 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(15, 5) & to_unsigned(4555, 13) & to_unsigned(4410, 13) & (12 downto 0 => 'U')),
    76 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(16, 5) & to_unsigned(4925, 13) & to_unsigned(4842, 13) & (12 downto 0 => 'U')),
    77 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(17, 5) & to_unsigned(5778, 13) & to_unsigned(600, 13) & (12 downto 0 => 'U')),
    78 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(18, 5) & to_unsigned(6509, 13) & to_unsigned(2417, 13) & (12 downto 0 => 'U')),
    79 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(19, 5) & to_unsigned(1260, 13) & to_unsigned(4903, 13) & (12 downto 0 => 'U')),
    80 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 5) & to_unsigned(3369, 13) & to_unsigned(3031, 13) & (12 downto 0 => 'U')),
    81 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 5) & to_unsigned(3557, 13) & to_unsigned(3224, 13) & (12 downto 0 => 'U')),
    82 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 5) & to_unsigned(3028, 13) & to_unsigned(583, 13) & (12 downto 0 => 'U')),
    83 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 5) & to_unsigned(3258, 13) & to_unsigned(440, 13) & (12 downto 0 => 'U')),
    84 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 5) & to_unsigned(6226, 13) & to_unsigned(6655, 13) & (12 downto 0 => 'U')),
    85 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(5, 5) & to_unsigned(4895, 13) & to_unsigned(1094, 13) & (12 downto 0 => 'U')),
    86 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(6, 5) & to_unsigned(1481, 13) & to_unsigned(6847, 13) & (12 downto 0 => 'U')),
    87 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(7, 5) & to_unsigned(4433, 13) & to_unsigned(1932, 13) & (12 downto 0 => 'U')),
    88 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(8, 5) & to_unsigned(2107, 13) & to_unsigned(1649, 13) & (12 downto 0 => 'U')),
    89 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(9, 5) & to_unsigned(2119, 13) & to_unsigned(2065, 13) & (12 downto 0 => 'U')),
    90 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(10, 5) & to_unsigned(4003, 13) & to_unsigned(6388, 13) & (12 downto 0 => 'U')),
    91 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(11, 5) & to_unsigned(6720, 13) & to_unsigned(3622, 13) & (12 downto 0 => 'U')),
    92 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(12, 5) & to_unsigned(3694, 13) & to_unsigned(4521, 13) & (12 downto 0 => 'U')),
    93 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(13, 5) & to_unsigned(1164, 13) & to_unsigned(7050, 13) & (12 downto 0 => 'U')),
    94 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(14, 5) & to_unsigned(1965, 13) & to_unsigned(3613, 13) & (12 downto 0 => 'U')),
    95 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(15, 5) & to_unsigned(4331, 13) & to_unsigned(66, 13) & (12 downto 0 => 'U')),
    96 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(16, 5) & to_unsigned(2970, 13) & to_unsigned(1796, 13) & (12 downto 0 => 'U')),
    97 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(17, 5) & to_unsigned(4652, 13) & to_unsigned(3218, 13) & (12 downto 0 => 'U')),
    98 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(18, 5) & to_unsigned(1762, 13) & to_unsigned(4777, 13) & (12 downto 0 => 'U')),
    99 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(19, 5) & to_unsigned(5736, 13) & to_unsigned(1399, 13) & (12 downto 0 => 'U')),
    100 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 5) & to_unsigned(970, 13) & to_unsigned(2572, 13) & (12 downto 0 => 'U')),
    101 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 5) & to_unsigned(2062, 13) & to_unsigned(6599, 13) & (12 downto 0 => 'U')),
    102 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 5) & to_unsigned(4597, 13) & to_unsigned(4870, 13) & (12 downto 0 => 'U')),
    103 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 5) & to_unsigned(1228, 13) & to_unsigned(6913, 13) & (12 downto 0 => 'U')),
    104 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 5) & to_unsigned(4159, 13) & to_unsigned(1037, 13) & (12 downto 0 => 'U')),
    105 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(5, 5) & to_unsigned(2916, 13) & to_unsigned(2362, 13) & (12 downto 0 => 'U')),
    106 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(6, 5) & to_unsigned(395, 13) & to_unsigned(1226, 13) & (12 downto 0 => 'U')),
    107 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(7, 5) & to_unsigned(6911, 13) & to_unsigned(4548, 13) & (12 downto 0 => 'U')),
    108 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(8, 5) & to_unsigned(4618, 13) & to_unsigned(2241, 13) & (12 downto 0 => 'U')),
    109 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(9, 5) & to_unsigned(4120, 13) & to_unsigned(4280, 13) & (12 downto 0 => 'U')),
    110 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(10, 5) & to_unsigned(5825, 13) & to_unsigned(474, 13) & (12 downto 0 => 'U')),
    111 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(11, 5) & to_unsigned(2154, 13) & to_unsigned(5558, 13) & (12 downto 0 => 'U')),
    112 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(12, 5) & to_unsigned(3793, 13) & to_unsigned(5471, 13) & (12 downto 0 => 'U')),
    113 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(13, 5) & to_unsigned(5707, 13) & to_unsigned(1595, 13) & (12 downto 0 => 'U')),
    114 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(14, 5) & to_unsigned(1403, 13) & to_unsigned(325, 13) & (12 downto 0 => 'U')),
    115 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(15, 5) & to_unsigned(6601, 13) & to_unsigned(5183, 13) & (12 downto 0 => 'U')),
    116 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(16, 5) & to_unsigned(6369, 13) & to_unsigned(4569, 13) & (12 downto 0 => 'U')),
    117 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(17, 5) & to_unsigned(4846, 13) & to_unsigned(896, 13) & (12 downto 0 => 'U')),
    118 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(18, 5) & to_unsigned(7092, 13) & to_unsigned(6184, 13) & (12 downto 0 => 'U')),
    119 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(19, 5) & to_unsigned(6764, 13) & to_unsigned(7127, 13) & (12 downto 0 => 'U')),
    120 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 5) & to_unsigned(6358, 13) & to_unsigned(1951, 13) & (12 downto 0 => 'U')),
    121 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 5) & to_unsigned(3117, 13) & to_unsigned(6960, 13) & (12 downto 0 => 'U')),
    122 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 5) & to_unsigned(2710, 13) & to_unsigned(7062, 13) & (12 downto 0 => 'U')),
    123 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 5) & to_unsigned(1133, 13) & to_unsigned(3604, 13) & (12 downto 0 => 'U')),
    124 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 5) & to_unsigned(3694, 13) & to_unsigned(657, 13) & (12 downto 0 => 'U')),
    125 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(5, 5) & to_unsigned(1355, 13) & to_unsigned(110, 13) & (12 downto 0 => 'U')),
    126 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(6, 5) & to_unsigned(3329, 13) & to_unsigned(6736, 13) & (12 downto 0 => 'U')),
    127 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(7, 5) & to_unsigned(2505, 13) & to_unsigned(3407, 13) & (12 downto 0 => 'U')),
    128 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(8, 5) & to_unsigned(2462, 13) & to_unsigned(4806, 13) & (12 downto 0 => 'U')),
    129 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(9, 5) & to_unsigned(4216, 13) & to_unsigned(214, 13) & (12 downto 0 => 'U')),
    130 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(10, 5) & to_unsigned(5348, 13) & to_unsigned(5619, 13) & (12 downto 0 => 'U')),
    131 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(11, 5) & to_unsigned(6627, 13) & to_unsigned(6243, 13) & (12 downto 0 => 'U')),
    132 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(12, 5) & to_unsigned(2644, 13) & to_unsigned(5073, 13) & (12 downto 0 => 'U')),
    133 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(13, 5) & to_unsigned(4212, 13) & to_unsigned(5088, 13) & (12 downto 0 => 'U')),
    134 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(14, 5) & to_unsigned(3463, 13) & to_unsigned(3889, 13) & (12 downto 0 => 'U')),
    135 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(15, 5) & to_unsigned(5306, 13) & to_unsigned(478, 13) & (12 downto 0 => 'U')),
    136 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(16, 5) & to_unsigned(4320, 13) & to_unsigned(6121, 13) & (12 downto 0 => 'U')),
    137 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(17, 5) & to_unsigned(3961, 13) & to_unsigned(1125, 13) & (12 downto 0 => 'U')),
    138 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(18, 5) & to_unsigned(5699, 13) & to_unsigned(1195, 13) & (12 downto 0 => 'U')),
    139 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(19, 5) & to_unsigned(6511, 13) & to_unsigned(792, 13) & (12 downto 0 => 'U')),
    140 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 5) & to_unsigned(3934, 13) & to_unsigned(2778, 13) & (12 downto 0 => 'U')),
    141 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 5) & to_unsigned(3238, 13) & to_unsigned(6587, 13) & (12 downto 0 => 'U')),
    142 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 5) & to_unsigned(1111, 13) & to_unsigned(6596, 13) & (12 downto 0 => 'U')),
    143 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 5) & to_unsigned(1457, 13) & to_unsigned(6226, 13) & (12 downto 0 => 'U')),
    144 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 5) & to_unsigned(1446, 13) & to_unsigned(3885, 13) & (12 downto 0 => 'U')),
    145 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(5, 5) & to_unsigned(3907, 13) & to_unsigned(4043, 13) & (12 downto 0 => 'U')),
    146 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(6, 5) & to_unsigned(6839, 13) & to_unsigned(2873, 13) & (12 downto 0 => 'U')),
    147 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(7, 5) & to_unsigned(1733, 13) & to_unsigned(5615, 13) & (12 downto 0 => 'U')),
    148 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(8, 5) & to_unsigned(5202, 13) & to_unsigned(4269, 13) & (12 downto 0 => 'U')),
    149 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(9, 5) & to_unsigned(3024, 13) & to_unsigned(4722, 13) & (12 downto 0 => 'U')),
    150 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(10, 5) & to_unsigned(5445, 13) & to_unsigned(6372, 13) & (12 downto 0 => 'U')),
    151 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(11, 5) & to_unsigned(370, 13) & to_unsigned(1828, 13) & (12 downto 0 => 'U')),
    152 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(12, 5) & to_unsigned(4695, 13) & to_unsigned(1600, 13) & (12 downto 0 => 'U')),
    153 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(13, 5) & to_unsigned(680, 13) & to_unsigned(2074, 13) & (12 downto 0 => 'U')),
    154 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(14, 5) & to_unsigned(1801, 13) & to_unsigned(6690, 13) & (12 downto 0 => 'U')),
    155 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(15, 5) & to_unsigned(2669, 13) & to_unsigned(1377, 13) & (12 downto 0 => 'U')),
    156 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(16, 5) & to_unsigned(2463, 13) & to_unsigned(1681, 13) & (12 downto 0 => 'U')),
    157 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(17, 5) & to_unsigned(5972, 13) & to_unsigned(5171, 13) & (12 downto 0 => 'U')),
    158 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(18, 5) & to_unsigned(5728, 13) & to_unsigned(4284, 13) & (12 downto 0 => 'U')),
    159 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(19, 5) & to_unsigned(1696, 13) & to_unsigned(1459, 13) & (12 downto 0 => 'U'))
  );

  -- From /home/souto/phase4ground/tables/ldpc/dvb/orig/dvb_64800_s2_b11.txt, table is 162x46 (931.5 bytes)
  -- Resource estimation: 3 x 18 kB BRAMs or 2 x 36 kB BRAMs
  type dvb_64800_s2_b11_t is array (161 downto 0) of std_logic_vector(45 downto 0);

  constant DVB_64800_S2_B11_COLUMN_WIDTHS : integer_array_t := (0 => 2, 1 => 5, 2 => 13, 3 => 13, 4 => 13);

  constant DVB_64800_S2_B11 : dvb_64800_s2_b11_t := (
    0 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(0, 5) & to_unsigned(5611, 13) & to_unsigned(2563, 13) & to_unsigned(2900, 13)),
    1 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(1, 5) & to_unsigned(5220, 13) & to_unsigned(3143, 13) & to_unsigned(4813, 13)),
    2 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(2, 5) & to_unsigned(2481, 13) & to_unsigned(834, 13) & to_unsigned(81, 13)),
    3 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(3, 5) & to_unsigned(6265, 13) & to_unsigned(4064, 13) & to_unsigned(4265, 13)),
    4 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(4, 5) & to_unsigned(1055, 13) & to_unsigned(2914, 13) & to_unsigned(5638, 13)),
    5 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(5, 5) & to_unsigned(1734, 13) & to_unsigned(2182, 13) & to_unsigned(3315, 13)),
    6 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(6, 5) & to_unsigned(3342, 13) & to_unsigned(5678, 13) & to_unsigned(2246, 13)),
    7 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(7, 5) & to_unsigned(2185, 13) & to_unsigned(552, 13) & to_unsigned(3385, 13)),
    8 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(8, 5) & to_unsigned(2615, 13) & to_unsigned(236, 13) & to_unsigned(5334, 13)),
    9 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(9, 5) & to_unsigned(1546, 13) & to_unsigned(1755, 13) & to_unsigned(3846, 13)),
    10 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(10, 5) & to_unsigned(4154, 13) & to_unsigned(5561, 13) & to_unsigned(3142, 13)),
    11 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(11, 5) & to_unsigned(4382, 13) & to_unsigned(2957, 13) & to_unsigned(5400, 13)),
    12 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(12, 5) & to_unsigned(1209, 13) & to_unsigned(5329, 13) & to_unsigned(3179, 13)),
    13 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(13, 5) & to_unsigned(1421, 13) & to_unsigned(3528, 13) & to_unsigned(6063, 13)),
    14 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(14, 5) & to_unsigned(1480, 13) & to_unsigned(1072, 13) & to_unsigned(5398, 13)),
    15 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(15, 5) & to_unsigned(3843, 13) & to_unsigned(1777, 13) & to_unsigned(4369, 13)),
    16 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(16, 5) & to_unsigned(1334, 13) & to_unsigned(2145, 13) & to_unsigned(4163, 13)),
    17 => std_logic_vector(to_unsigned(4, 2) & to_unsigned(17, 5) & to_unsigned(2368, 13) & to_unsigned(5055, 13) & to_unsigned(260, 13)),
    18 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 5) & to_unsigned(6118, 13) & to_unsigned(5405, 13) & (12 downto 0 => 'U')),
    19 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 5) & to_unsigned(2994, 13) & to_unsigned(4370, 13) & (12 downto 0 => 'U')),
    20 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 5) & to_unsigned(3405, 13) & to_unsigned(1669, 13) & (12 downto 0 => 'U')),
    21 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 5) & to_unsigned(4640, 13) & to_unsigned(5550, 13) & (12 downto 0 => 'U')),
    22 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 5) & to_unsigned(1354, 13) & to_unsigned(3921, 13) & (12 downto 0 => 'U')),
    23 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(5, 5) & to_unsigned(117, 13) & to_unsigned(1713, 13) & (12 downto 0 => 'U')),
    24 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(6, 5) & to_unsigned(5425, 13) & to_unsigned(2866, 13) & (12 downto 0 => 'U')),
    25 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(7, 5) & to_unsigned(6047, 13) & to_unsigned(683, 13) & (12 downto 0 => 'U')),
    26 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(8, 5) & to_unsigned(5616, 13) & to_unsigned(2582, 13) & (12 downto 0 => 'U')),
    27 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(9, 5) & to_unsigned(2108, 13) & to_unsigned(1179, 13) & (12 downto 0 => 'U')),
    28 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(10, 5) & to_unsigned(933, 13) & to_unsigned(4921, 13) & (12 downto 0 => 'U')),
    29 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(11, 5) & to_unsigned(5953, 13) & to_unsigned(2261, 13) & (12 downto 0 => 'U')),
    30 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(12, 5) & to_unsigned(1430, 13) & to_unsigned(4699, 13) & (12 downto 0 => 'U')),
    31 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(13, 5) & to_unsigned(5905, 13) & to_unsigned(480, 13) & (12 downto 0 => 'U')),
    32 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(14, 5) & to_unsigned(4289, 13) & to_unsigned(1846, 13) & (12 downto 0 => 'U')),
    33 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(15, 5) & to_unsigned(5374, 13) & to_unsigned(6208, 13) & (12 downto 0 => 'U')),
    34 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(16, 5) & to_unsigned(1775, 13) & to_unsigned(3476, 13) & (12 downto 0 => 'U')),
    35 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(17, 5) & to_unsigned(3216, 13) & to_unsigned(2178, 13) & (12 downto 0 => 'U')),
    36 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 5) & to_unsigned(4165, 13) & to_unsigned(884, 13) & (12 downto 0 => 'U')),
    37 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 5) & to_unsigned(2896, 13) & to_unsigned(3744, 13) & (12 downto 0 => 'U')),
    38 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 5) & to_unsigned(874, 13) & to_unsigned(2801, 13) & (12 downto 0 => 'U')),
    39 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 5) & to_unsigned(3423, 13) & to_unsigned(5579, 13) & (12 downto 0 => 'U')),
    40 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 5) & to_unsigned(3404, 13) & to_unsigned(3552, 13) & (12 downto 0 => 'U')),
    41 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(5, 5) & to_unsigned(2876, 13) & to_unsigned(5515, 13) & (12 downto 0 => 'U')),
    42 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(6, 5) & to_unsigned(516, 13) & to_unsigned(1719, 13) & (12 downto 0 => 'U')),
    43 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(7, 5) & to_unsigned(765, 13) & to_unsigned(3631, 13) & (12 downto 0 => 'U')),
    44 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(8, 5) & to_unsigned(5059, 13) & to_unsigned(1441, 13) & (12 downto 0 => 'U')),
    45 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(9, 5) & to_unsigned(5629, 13) & to_unsigned(598, 13) & (12 downto 0 => 'U')),
    46 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(10, 5) & to_unsigned(5405, 13) & to_unsigned(473, 13) & (12 downto 0 => 'U')),
    47 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(11, 5) & to_unsigned(4724, 13) & to_unsigned(5210, 13) & (12 downto 0 => 'U')),
    48 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(12, 5) & to_unsigned(155, 13) & to_unsigned(1832, 13) & (12 downto 0 => 'U')),
    49 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(13, 5) & to_unsigned(1689, 13) & to_unsigned(2229, 13) & (12 downto 0 => 'U')),
    50 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(14, 5) & to_unsigned(449, 13) & to_unsigned(1164, 13) & (12 downto 0 => 'U')),
    51 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(15, 5) & to_unsigned(2308, 13) & to_unsigned(3088, 13) & (12 downto 0 => 'U')),
    52 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(16, 5) & to_unsigned(1122, 13) & to_unsigned(669, 13) & (12 downto 0 => 'U')),
    53 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(17, 5) & to_unsigned(2268, 13) & to_unsigned(5758, 13) & (12 downto 0 => 'U')),
    54 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 5) & to_unsigned(5878, 13) & to_unsigned(2609, 13) & (12 downto 0 => 'U')),
    55 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 5) & to_unsigned(782, 13) & to_unsigned(3359, 13) & (12 downto 0 => 'U')),
    56 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 5) & to_unsigned(1231, 13) & to_unsigned(4231, 13) & (12 downto 0 => 'U')),
    57 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 5) & to_unsigned(4225, 13) & to_unsigned(2052, 13) & (12 downto 0 => 'U')),
    58 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 5) & to_unsigned(4286, 13) & to_unsigned(3517, 13) & (12 downto 0 => 'U')),
    59 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(5, 5) & to_unsigned(5531, 13) & to_unsigned(3184, 13) & (12 downto 0 => 'U')),
    60 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(6, 5) & to_unsigned(1935, 13) & to_unsigned(4560, 13) & (12 downto 0 => 'U')),
    61 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(7, 5) & to_unsigned(1174, 13) & to_unsigned(131, 13) & (12 downto 0 => 'U')),
    62 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(8, 5) & to_unsigned(3115, 13) & to_unsigned(956, 13) & (12 downto 0 => 'U')),
    63 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(9, 5) & to_unsigned(3129, 13) & to_unsigned(1088, 13) & (12 downto 0 => 'U')),
    64 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(10, 5) & to_unsigned(5238, 13) & to_unsigned(4440, 13) & (12 downto 0 => 'U')),
    65 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(11, 5) & to_unsigned(5722, 13) & to_unsigned(4280, 13) & (12 downto 0 => 'U')),
    66 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(12, 5) & to_unsigned(3540, 13) & to_unsigned(375, 13) & (12 downto 0 => 'U')),
    67 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(13, 5) & to_unsigned(191, 13) & to_unsigned(2782, 13) & (12 downto 0 => 'U')),
    68 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(14, 5) & to_unsigned(906, 13) & to_unsigned(4432, 13) & (12 downto 0 => 'U')),
    69 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(15, 5) & to_unsigned(3225, 13) & to_unsigned(1111, 13) & (12 downto 0 => 'U')),
    70 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(16, 5) & to_unsigned(6296, 13) & to_unsigned(2583, 13) & (12 downto 0 => 'U')),
    71 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(17, 5) & to_unsigned(1457, 13) & to_unsigned(903, 13) & (12 downto 0 => 'U')),
    72 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 5) & to_unsigned(855, 13) & to_unsigned(4475, 13) & (12 downto 0 => 'U')),
    73 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 5) & to_unsigned(4097, 13) & to_unsigned(3970, 13) & (12 downto 0 => 'U')),
    74 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 5) & to_unsigned(4433, 13) & to_unsigned(4361, 13) & (12 downto 0 => 'U')),
    75 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 5) & to_unsigned(5198, 13) & to_unsigned(541, 13) & (12 downto 0 => 'U')),
    76 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 5) & to_unsigned(1146, 13) & to_unsigned(4426, 13) & (12 downto 0 => 'U')),
    77 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(5, 5) & to_unsigned(3202, 13) & to_unsigned(2902, 13) & (12 downto 0 => 'U')),
    78 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(6, 5) & to_unsigned(2724, 13) & to_unsigned(525, 13) & (12 downto 0 => 'U')),
    79 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(7, 5) & to_unsigned(1083, 13) & to_unsigned(4124, 13) & (12 downto 0 => 'U')),
    80 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(8, 5) & to_unsigned(2326, 13) & to_unsigned(6003, 13) & (12 downto 0 => 'U')),
    81 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(9, 5) & to_unsigned(5605, 13) & to_unsigned(5990, 13) & (12 downto 0 => 'U')),
    82 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(10, 5) & to_unsigned(4376, 13) & to_unsigned(1579, 13) & (12 downto 0 => 'U')),
    83 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(11, 5) & to_unsigned(4407, 13) & to_unsigned(984, 13) & (12 downto 0 => 'U')),
    84 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(12, 5) & to_unsigned(1332, 13) & to_unsigned(6163, 13) & (12 downto 0 => 'U')),
    85 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(13, 5) & to_unsigned(5359, 13) & to_unsigned(3975, 13) & (12 downto 0 => 'U')),
    86 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(14, 5) & to_unsigned(1907, 13) & to_unsigned(1854, 13) & (12 downto 0 => 'U')),
    87 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(15, 5) & to_unsigned(3601, 13) & to_unsigned(5748, 13) & (12 downto 0 => 'U')),
    88 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(16, 5) & to_unsigned(6056, 13) & to_unsigned(3266, 13) & (12 downto 0 => 'U')),
    89 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(17, 5) & to_unsigned(3322, 13) & to_unsigned(4085, 13) & (12 downto 0 => 'U')),
    90 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 5) & to_unsigned(1768, 13) & to_unsigned(3244, 13) & (12 downto 0 => 'U')),
    91 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 5) & to_unsigned(2149, 13) & to_unsigned(144, 13) & (12 downto 0 => 'U')),
    92 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 5) & to_unsigned(1589, 13) & to_unsigned(4291, 13) & (12 downto 0 => 'U')),
    93 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 5) & to_unsigned(5154, 13) & to_unsigned(1252, 13) & (12 downto 0 => 'U')),
    94 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 5) & to_unsigned(1855, 13) & to_unsigned(5939, 13) & (12 downto 0 => 'U')),
    95 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(5, 5) & to_unsigned(4820, 13) & to_unsigned(2706, 13) & (12 downto 0 => 'U')),
    96 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(6, 5) & to_unsigned(1475, 13) & to_unsigned(3360, 13) & (12 downto 0 => 'U')),
    97 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(7, 5) & to_unsigned(4266, 13) & to_unsigned(693, 13) & (12 downto 0 => 'U')),
    98 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(8, 5) & to_unsigned(4156, 13) & to_unsigned(2018, 13) & (12 downto 0 => 'U')),
    99 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(9, 5) & to_unsigned(2103, 13) & to_unsigned(752, 13) & (12 downto 0 => 'U')),
    100 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(10, 5) & to_unsigned(3710, 13) & to_unsigned(3853, 13) & (12 downto 0 => 'U')),
    101 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(11, 5) & to_unsigned(5123, 13) & to_unsigned(931, 13) & (12 downto 0 => 'U')),
    102 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(12, 5) & to_unsigned(6146, 13) & to_unsigned(3323, 13) & (12 downto 0 => 'U')),
    103 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(13, 5) & to_unsigned(1939, 13) & to_unsigned(5002, 13) & (12 downto 0 => 'U')),
    104 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(14, 5) & to_unsigned(5140, 13) & to_unsigned(1437, 13) & (12 downto 0 => 'U')),
    105 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(15, 5) & to_unsigned(1263, 13) & to_unsigned(293, 13) & (12 downto 0 => 'U')),
    106 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(16, 5) & to_unsigned(5949, 13) & to_unsigned(4665, 13) & (12 downto 0 => 'U')),
    107 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(17, 5) & to_unsigned(4548, 13) & to_unsigned(6380, 13) & (12 downto 0 => 'U')),
    108 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 5) & to_unsigned(3171, 13) & to_unsigned(4690, 13) & (12 downto 0 => 'U')),
    109 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 5) & to_unsigned(5204, 13) & to_unsigned(2114, 13) & (12 downto 0 => 'U')),
    110 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 5) & to_unsigned(6384, 13) & to_unsigned(5565, 13) & (12 downto 0 => 'U')),
    111 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 5) & to_unsigned(5722, 13) & to_unsigned(1757, 13) & (12 downto 0 => 'U')),
    112 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 5) & to_unsigned(2805, 13) & to_unsigned(6264, 13) & (12 downto 0 => 'U')),
    113 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(5, 5) & to_unsigned(1202, 13) & to_unsigned(2616, 13) & (12 downto 0 => 'U')),
    114 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(6, 5) & to_unsigned(1018, 13) & to_unsigned(3244, 13) & (12 downto 0 => 'U')),
    115 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(7, 5) & to_unsigned(4018, 13) & to_unsigned(5289, 13) & (12 downto 0 => 'U')),
    116 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(8, 5) & to_unsigned(2257, 13) & to_unsigned(3067, 13) & (12 downto 0 => 'U')),
    117 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(9, 5) & to_unsigned(2483, 13) & to_unsigned(3073, 13) & (12 downto 0 => 'U')),
    118 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(10, 5) & to_unsigned(1196, 13) & to_unsigned(5329, 13) & (12 downto 0 => 'U')),
    119 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(11, 5) & to_unsigned(649, 13) & to_unsigned(3918, 13) & (12 downto 0 => 'U')),
    120 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(12, 5) & to_unsigned(3791, 13) & to_unsigned(4581, 13) & (12 downto 0 => 'U')),
    121 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(13, 5) & to_unsigned(5028, 13) & to_unsigned(3803, 13) & (12 downto 0 => 'U')),
    122 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(14, 5) & to_unsigned(3119, 13) & to_unsigned(3506, 13) & (12 downto 0 => 'U')),
    123 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(15, 5) & to_unsigned(4779, 13) & to_unsigned(431, 13) & (12 downto 0 => 'U')),
    124 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(16, 5) & to_unsigned(3888, 13) & to_unsigned(5510, 13) & (12 downto 0 => 'U')),
    125 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(17, 5) & to_unsigned(4387, 13) & to_unsigned(4084, 13) & (12 downto 0 => 'U')),
    126 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 5) & to_unsigned(5836, 13) & to_unsigned(1692, 13) & (12 downto 0 => 'U')),
    127 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 5) & to_unsigned(5126, 13) & to_unsigned(1078, 13) & (12 downto 0 => 'U')),
    128 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 5) & to_unsigned(5721, 13) & to_unsigned(6165, 13) & (12 downto 0 => 'U')),
    129 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 5) & to_unsigned(3540, 13) & to_unsigned(2499, 13) & (12 downto 0 => 'U')),
    130 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 5) & to_unsigned(2225, 13) & to_unsigned(6348, 13) & (12 downto 0 => 'U')),
    131 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(5, 5) & to_unsigned(1044, 13) & to_unsigned(1484, 13) & (12 downto 0 => 'U')),
    132 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(6, 5) & to_unsigned(6323, 13) & to_unsigned(4042, 13) & (12 downto 0 => 'U')),
    133 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(7, 5) & to_unsigned(1313, 13) & to_unsigned(5603, 13) & (12 downto 0 => 'U')),
    134 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(8, 5) & to_unsigned(1303, 13) & to_unsigned(3496, 13) & (12 downto 0 => 'U')),
    135 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(9, 5) & to_unsigned(3516, 13) & to_unsigned(3639, 13) & (12 downto 0 => 'U')),
    136 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(10, 5) & to_unsigned(5161, 13) & to_unsigned(2293, 13) & (12 downto 0 => 'U')),
    137 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(11, 5) & to_unsigned(4682, 13) & to_unsigned(3845, 13) & (12 downto 0 => 'U')),
    138 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(12, 5) & to_unsigned(3045, 13) & to_unsigned(643, 13) & (12 downto 0 => 'U')),
    139 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(13, 5) & to_unsigned(2818, 13) & to_unsigned(2616, 13) & (12 downto 0 => 'U')),
    140 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(14, 5) & to_unsigned(3267, 13) & to_unsigned(649, 13) & (12 downto 0 => 'U')),
    141 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(15, 5) & to_unsigned(6236, 13) & to_unsigned(593, 13) & (12 downto 0 => 'U')),
    142 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(16, 5) & to_unsigned(646, 13) & to_unsigned(2948, 13) & (12 downto 0 => 'U')),
    143 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(17, 5) & to_unsigned(4213, 13) & to_unsigned(1442, 13) & (12 downto 0 => 'U')),
    144 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(0, 5) & to_unsigned(5779, 13) & to_unsigned(1596, 13) & (12 downto 0 => 'U')),
    145 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(1, 5) & to_unsigned(2403, 13) & to_unsigned(1237, 13) & (12 downto 0 => 'U')),
    146 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(2, 5) & to_unsigned(2217, 13) & to_unsigned(1514, 13) & (12 downto 0 => 'U')),
    147 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(3, 5) & to_unsigned(5609, 13) & to_unsigned(716, 13) & (12 downto 0 => 'U')),
    148 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(4, 5) & to_unsigned(5155, 13) & to_unsigned(3858, 13) & (12 downto 0 => 'U')),
    149 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(5, 5) & to_unsigned(1517, 13) & to_unsigned(1312, 13) & (12 downto 0 => 'U')),
    150 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(6, 5) & to_unsigned(2554, 13) & to_unsigned(3158, 13) & (12 downto 0 => 'U')),
    151 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(7, 5) & to_unsigned(5280, 13) & to_unsigned(2643, 13) & (12 downto 0 => 'U')),
    152 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(8, 5) & to_unsigned(4990, 13) & to_unsigned(1353, 13) & (12 downto 0 => 'U')),
    153 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(9, 5) & to_unsigned(5648, 13) & to_unsigned(1170, 13) & (12 downto 0 => 'U')),
    154 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(10, 5) & to_unsigned(1152, 13) & to_unsigned(4366, 13) & (12 downto 0 => 'U')),
    155 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(11, 5) & to_unsigned(3561, 13) & to_unsigned(5368, 13) & (12 downto 0 => 'U')),
    156 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(12, 5) & to_unsigned(3581, 13) & to_unsigned(1411, 13) & (12 downto 0 => 'U')),
    157 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(13, 5) & to_unsigned(5647, 13) & to_unsigned(4661, 13) & (12 downto 0 => 'U')),
    158 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(14, 5) & to_unsigned(1542, 13) & to_unsigned(5401, 13) & (12 downto 0 => 'U')),
    159 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(15, 5) & to_unsigned(5078, 13) & to_unsigned(2687, 13) & (12 downto 0 => 'U')),
    160 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(16, 5) & to_unsigned(316, 13) & to_unsigned(1755, 13) & (12 downto 0 => 'U')),
    161 => std_logic_vector(to_unsigned(3, 2) & to_unsigned(17, 5) & to_unsigned(3392, 13) & to_unsigned(1991, 13) & (12 downto 0 => 'U'))
  );

  -- From /home/souto/phase4ground/tables/ldpc/dvb/orig/dvb_64800_s2_b2.txt, table is 60x196 (1470.0 bytes)
  -- Resource estimation: 11 x 18 kB BRAMs or 6 x 36 kB BRAMs
  type dvb_64800_s2_b2_t is array (59 downto 0) of std_logic_vector(195 downto 0);

  constant DVB_64800_S2_B2_COLUMN_WIDTHS : integer_array_t := (0 => 4, 1 => 16, 2 => 16, 3 => 16, 4 => 16, 5 => 16, 6 => 16, 7 => 16, 8 => 16, 9 => 16, 10 => 16, 11 => 16, 12 => 16);

  constant DVB_64800_S2_B2 : dvb_64800_s2_b2_t := (
    0 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(34903, 16) & to_unsigned(20927, 16) & to_unsigned(32093, 16) & to_unsigned(1052, 16) & to_unsigned(25611, 16) & to_unsigned(16093, 16) & to_unsigned(16454, 16) & to_unsigned(5520, 16) & to_unsigned(506, 16) & to_unsigned(37399, 16) & to_unsigned(18518, 16) & to_unsigned(21120, 16)),
    1 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(11636, 16) & to_unsigned(14594, 16) & to_unsigned(22158, 16) & to_unsigned(14763, 16) & to_unsigned(15333, 16) & to_unsigned(6838, 16) & to_unsigned(22222, 16) & to_unsigned(37856, 16) & to_unsigned(14985, 16) & to_unsigned(31041, 16) & to_unsigned(18704, 16) & to_unsigned(32910, 16)),
    2 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(17449, 16) & to_unsigned(1665, 16) & to_unsigned(35639, 16) & to_unsigned(16624, 16) & to_unsigned(12867, 16) & to_unsigned(12449, 16) & to_unsigned(10241, 16) & to_unsigned(11650, 16) & to_unsigned(25622, 16) & to_unsigned(34372, 16) & to_unsigned(19878, 16) & to_unsigned(26894, 16)),
    3 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(29235, 16) & to_unsigned(19780, 16) & to_unsigned(36056, 16) & to_unsigned(20129, 16) & to_unsigned(20029, 16) & to_unsigned(5457, 16) & to_unsigned(8157, 16) & to_unsigned(35554, 16) & to_unsigned(21237, 16) & to_unsigned(7943, 16) & to_unsigned(13873, 16) & to_unsigned(14980, 16)),
    4 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(9912, 16) & to_unsigned(7143, 16) & to_unsigned(35911, 16) & to_unsigned(12043, 16) & to_unsigned(17360, 16) & to_unsigned(37253, 16) & to_unsigned(25588, 16) & to_unsigned(11827, 16) & to_unsigned(29152, 16) & to_unsigned(21936, 16) & to_unsigned(24125, 16) & to_unsigned(40870, 16)),
    5 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(40701, 16) & to_unsigned(36035, 16) & to_unsigned(39556, 16) & to_unsigned(12366, 16) & to_unsigned(19946, 16) & to_unsigned(29072, 16) & to_unsigned(16365, 16) & to_unsigned(35495, 16) & to_unsigned(22686, 16) & to_unsigned(11106, 16) & to_unsigned(8756, 16) & to_unsigned(34863, 16)),
    6 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(19165, 16) & to_unsigned(15702, 16) & to_unsigned(13536, 16) & to_unsigned(40238, 16) & to_unsigned(4465, 16) & to_unsigned(40034, 16) & to_unsigned(40590, 16) & to_unsigned(37540, 16) & to_unsigned(17162, 16) & to_unsigned(1712, 16) & to_unsigned(20577, 16) & to_unsigned(14138, 16)),
    7 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(31338, 16) & to_unsigned(19342, 16) & to_unsigned(9301, 16) & to_unsigned(39375, 16) & to_unsigned(3211, 16) & to_unsigned(1316, 16) & to_unsigned(33409, 16) & to_unsigned(28670, 16) & to_unsigned(12282, 16) & to_unsigned(6118, 16) & to_unsigned(29236, 16) & to_unsigned(35787, 16)),
    8 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(11504, 16) & to_unsigned(30506, 16) & to_unsigned(19558, 16) & to_unsigned(5100, 16) & to_unsigned(24188, 16) & to_unsigned(24738, 16) & to_unsigned(30397, 16) & to_unsigned(33775, 16) & to_unsigned(9699, 16) & to_unsigned(6215, 16) & to_unsigned(3397, 16) & to_unsigned(37451, 16)),
    9 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(34689, 16) & to_unsigned(23126, 16) & to_unsigned(7571, 16) & to_unsigned(1058, 16) & to_unsigned(12127, 16) & to_unsigned(27518, 16) & to_unsigned(23064, 16) & to_unsigned(11265, 16) & to_unsigned(14867, 16) & to_unsigned(30451, 16) & to_unsigned(28289, 16) & to_unsigned(2966, 16)),
    10 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(11660, 16) & to_unsigned(15334, 16) & to_unsigned(16867, 16) & to_unsigned(15160, 16) & to_unsigned(38343, 16) & to_unsigned(3778, 16) & to_unsigned(4265, 16) & to_unsigned(39139, 16) & to_unsigned(17293, 16) & to_unsigned(26229, 16) & to_unsigned(42604, 16) & to_unsigned(13486, 16)),
    11 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(31497, 16) & to_unsigned(1365, 16) & to_unsigned(14828, 16) & to_unsigned(7453, 16) & to_unsigned(26350, 16) & to_unsigned(41346, 16) & to_unsigned(28643, 16) & to_unsigned(23421, 16) & to_unsigned(8354, 16) & to_unsigned(16255, 16) & to_unsigned(11055, 16) & to_unsigned(24279, 16)),
    12 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(15687, 16) & to_unsigned(12467, 16) & to_unsigned(13906, 16) & to_unsigned(5215, 16) & to_unsigned(41328, 16) & to_unsigned(23755, 16) & to_unsigned(20800, 16) & to_unsigned(6447, 16) & to_unsigned(7970, 16) & to_unsigned(2803, 16) & to_unsigned(33262, 16) & to_unsigned(39843, 16)),
    13 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(5363, 16) & to_unsigned(22469, 16) & to_unsigned(38091, 16) & to_unsigned(28457, 16) & to_unsigned(36696, 16) & to_unsigned(34471, 16) & to_unsigned(23619, 16) & to_unsigned(2404, 16) & to_unsigned(24229, 16) & to_unsigned(41754, 16) & to_unsigned(1297, 16) & to_unsigned(18563, 16)),
    14 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(3673, 16) & to_unsigned(39070, 16) & to_unsigned(14480, 16) & to_unsigned(30279, 16) & to_unsigned(37483, 16) & to_unsigned(7580, 16) & to_unsigned(29519, 16) & to_unsigned(30519, 16) & to_unsigned(39831, 16) & to_unsigned(20252, 16) & to_unsigned(18132, 16) & to_unsigned(20010, 16)),
    15 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(34386, 16) & to_unsigned(7252, 16) & to_unsigned(27526, 16) & to_unsigned(12950, 16) & to_unsigned(6875, 16) & to_unsigned(43020, 16) & to_unsigned(31566, 16) & to_unsigned(39069, 16) & to_unsigned(18985, 16) & to_unsigned(15541, 16) & to_unsigned(40020, 16) & to_unsigned(16715, 16)),
    16 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(1721, 16) & to_unsigned(37332, 16) & to_unsigned(39953, 16) & to_unsigned(17430, 16) & to_unsigned(32134, 16) & to_unsigned(29162, 16) & to_unsigned(10490, 16) & to_unsigned(12971, 16) & to_unsigned(28581, 16) & to_unsigned(29331, 16) & to_unsigned(6489, 16) & to_unsigned(35383, 16)),
    17 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(736, 16) & to_unsigned(7022, 16) & to_unsigned(42349, 16) & to_unsigned(8783, 16) & to_unsigned(6767, 16) & to_unsigned(11871, 16) & to_unsigned(21675, 16) & to_unsigned(10325, 16) & to_unsigned(11548, 16) & to_unsigned(25978, 16) & to_unsigned(431, 16) & to_unsigned(24085, 16)),
    18 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(1925, 16) & to_unsigned(10602, 16) & to_unsigned(28585, 16) & to_unsigned(12170, 16) & to_unsigned(15156, 16) & to_unsigned(34404, 16) & to_unsigned(8351, 16) & to_unsigned(13273, 16) & to_unsigned(20208, 16) & to_unsigned(5800, 16) & to_unsigned(15367, 16) & to_unsigned(21764, 16)),
    19 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(16279, 16) & to_unsigned(37832, 16) & to_unsigned(34792, 16) & to_unsigned(21250, 16) & to_unsigned(34192, 16) & to_unsigned(7406, 16) & to_unsigned(41488, 16) & to_unsigned(18346, 16) & to_unsigned(29227, 16) & to_unsigned(26127, 16) & to_unsigned(25493, 16) & to_unsigned(7048, 16)),
    20 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(39948, 16) & to_unsigned(28229, 16) & to_unsigned(24899, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    21 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(17408, 16) & to_unsigned(14274, 16) & to_unsigned(38993, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    22 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(38774, 16) & to_unsigned(15968, 16) & to_unsigned(28459, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    23 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(41404, 16) & to_unsigned(27249, 16) & to_unsigned(27425, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    24 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(41229, 16) & to_unsigned(6082, 16) & to_unsigned(43114, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    25 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(13957, 16) & to_unsigned(4979, 16) & to_unsigned(40654, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    26 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3093, 16) & to_unsigned(3438, 16) & to_unsigned(34992, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    27 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(34082, 16) & to_unsigned(6172, 16) & to_unsigned(28760, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    28 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(42210, 16) & to_unsigned(34141, 16) & to_unsigned(41021, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    29 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(14705, 16) & to_unsigned(17783, 16) & to_unsigned(10134, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    30 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(41755, 16) & to_unsigned(39884, 16) & to_unsigned(22773, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    31 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(14615, 16) & to_unsigned(15593, 16) & to_unsigned(1642, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    32 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(29111, 16) & to_unsigned(37061, 16) & to_unsigned(39860, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    33 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9579, 16) & to_unsigned(33552, 16) & to_unsigned(633, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    34 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(12951, 16) & to_unsigned(21137, 16) & to_unsigned(39608, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    35 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(38244, 16) & to_unsigned(27361, 16) & to_unsigned(29417, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    36 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(2939, 16) & to_unsigned(10172, 16) & to_unsigned(36479, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    37 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(29094, 16) & to_unsigned(5357, 16) & to_unsigned(19224, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    38 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9562, 16) & to_unsigned(24436, 16) & to_unsigned(28637, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    39 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(40177, 16) & to_unsigned(2326, 16) & to_unsigned(13504, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    40 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6834, 16) & to_unsigned(21583, 16) & to_unsigned(42516, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    41 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(40651, 16) & to_unsigned(42810, 16) & to_unsigned(25709, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    42 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(31557, 16) & to_unsigned(32138, 16) & to_unsigned(38142, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    43 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(18624, 16) & to_unsigned(41867, 16) & to_unsigned(39296, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    44 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(37560, 16) & to_unsigned(14295, 16) & to_unsigned(16245, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    45 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6821, 16) & to_unsigned(21679, 16) & to_unsigned(31570, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    46 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(25339, 16) & to_unsigned(25083, 16) & to_unsigned(22081, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    47 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(8047, 16) & to_unsigned(697, 16) & to_unsigned(35268, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    48 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9884, 16) & to_unsigned(17073, 16) & to_unsigned(19995, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    49 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(26848, 16) & to_unsigned(35245, 16) & to_unsigned(8390, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    50 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(18658, 16) & to_unsigned(16134, 16) & to_unsigned(14807, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    51 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(12201, 16) & to_unsigned(32944, 16) & to_unsigned(5035, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    52 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(25236, 16) & to_unsigned(1216, 16) & to_unsigned(38986, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    53 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(42994, 16) & to_unsigned(24782, 16) & to_unsigned(8681, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    54 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(28321, 16) & to_unsigned(4932, 16) & to_unsigned(34249, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    55 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4107, 16) & to_unsigned(29382, 16) & to_unsigned(32124, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    56 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(22157, 16) & to_unsigned(2624, 16) & to_unsigned(14468, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    57 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(38788, 16) & to_unsigned(27081, 16) & to_unsigned(7936, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    58 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4368, 16) & to_unsigned(26148, 16) & to_unsigned(10578, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    59 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(25353, 16) & to_unsigned(4122, 16) & to_unsigned(39751, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U'))
  );

  -- From /home/souto/phase4ground/tables/ldpc/dvb/orig/dvb_64800_s2_b3.txt, table is 72x196 (1764.0 bytes)
  -- Resource estimation: 11 x 18 kB BRAMs or 6 x 36 kB BRAMs
  type dvb_64800_s2_b3_t is array (71 downto 0) of std_logic_vector(195 downto 0);

  constant DVB_64800_S2_B3_COLUMN_WIDTHS : integer_array_t := (0 => 4, 1 => 16, 2 => 16, 3 => 16, 4 => 16, 5 => 16, 6 => 16, 7 => 16, 8 => 16, 9 => 16, 10 => 16, 11 => 16, 12 => 16);

  constant DVB_64800_S2_B3 : dvb_64800_s2_b3_t := (
    0 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(31413, 16) & to_unsigned(18834, 16) & to_unsigned(28884, 16) & to_unsigned(947, 16) & to_unsigned(23050, 16) & to_unsigned(14484, 16) & to_unsigned(14809, 16) & to_unsigned(4968, 16) & to_unsigned(455, 16) & to_unsigned(33659, 16) & to_unsigned(16666, 16) & to_unsigned(19008, 16)),
    1 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(13172, 16) & to_unsigned(19939, 16) & to_unsigned(13354, 16) & to_unsigned(13719, 16) & to_unsigned(6132, 16) & to_unsigned(20086, 16) & to_unsigned(34040, 16) & to_unsigned(13442, 16) & to_unsigned(27958, 16) & to_unsigned(16813, 16) & to_unsigned(29619, 16) & to_unsigned(16553, 16)),
    2 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(1499, 16) & to_unsigned(32075, 16) & to_unsigned(14962, 16) & to_unsigned(11578, 16) & to_unsigned(11204, 16) & to_unsigned(9217, 16) & to_unsigned(10485, 16) & to_unsigned(23062, 16) & to_unsigned(30936, 16) & to_unsigned(17892, 16) & to_unsigned(24204, 16) & to_unsigned(24885, 16)),
    3 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(32490, 16) & to_unsigned(18086, 16) & to_unsigned(18007, 16) & to_unsigned(4957, 16) & to_unsigned(7285, 16) & to_unsigned(32073, 16) & to_unsigned(19038, 16) & to_unsigned(7152, 16) & to_unsigned(12486, 16) & to_unsigned(13483, 16) & to_unsigned(24808, 16) & to_unsigned(21759, 16)),
    4 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(32321, 16) & to_unsigned(10839, 16) & to_unsigned(15620, 16) & to_unsigned(33521, 16) & to_unsigned(23030, 16) & to_unsigned(10646, 16) & to_unsigned(26236, 16) & to_unsigned(19744, 16) & to_unsigned(21713, 16) & to_unsigned(36784, 16) & to_unsigned(8016, 16) & to_unsigned(12869, 16)),
    5 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(35597, 16) & to_unsigned(11129, 16) & to_unsigned(17948, 16) & to_unsigned(26160, 16) & to_unsigned(14729, 16) & to_unsigned(31943, 16) & to_unsigned(20416, 16) & to_unsigned(10000, 16) & to_unsigned(7882, 16) & to_unsigned(31380, 16) & to_unsigned(27858, 16) & to_unsigned(33356, 16)),
    6 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(14125, 16) & to_unsigned(12131, 16) & to_unsigned(36199, 16) & to_unsigned(4058, 16) & to_unsigned(35992, 16) & to_unsigned(36594, 16) & to_unsigned(33698, 16) & to_unsigned(15475, 16) & to_unsigned(1566, 16) & to_unsigned(18498, 16) & to_unsigned(12725, 16) & to_unsigned(7067, 16)),
    7 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(17406, 16) & to_unsigned(8372, 16) & to_unsigned(35437, 16) & to_unsigned(2888, 16) & to_unsigned(1184, 16) & to_unsigned(30068, 16) & to_unsigned(25802, 16) & to_unsigned(11056, 16) & to_unsigned(5507, 16) & to_unsigned(26313, 16) & to_unsigned(32205, 16) & to_unsigned(37232, 16)),
    8 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(15254, 16) & to_unsigned(5365, 16) & to_unsigned(17308, 16) & to_unsigned(22519, 16) & to_unsigned(35009, 16) & to_unsigned(718, 16) & to_unsigned(5240, 16) & to_unsigned(16778, 16) & to_unsigned(23131, 16) & to_unsigned(24092, 16) & to_unsigned(20587, 16) & to_unsigned(33385, 16)),
    9 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(27455, 16) & to_unsigned(17602, 16) & to_unsigned(4590, 16) & to_unsigned(21767, 16) & to_unsigned(22266, 16) & to_unsigned(27357, 16) & to_unsigned(30400, 16) & to_unsigned(8732, 16) & to_unsigned(5596, 16) & to_unsigned(3060, 16) & to_unsigned(33703, 16) & to_unsigned(3596, 16)),
    10 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(6882, 16) & to_unsigned(873, 16) & to_unsigned(10997, 16) & to_unsigned(24738, 16) & to_unsigned(20770, 16) & to_unsigned(10067, 16) & to_unsigned(13379, 16) & to_unsigned(27409, 16) & to_unsigned(25463, 16) & to_unsigned(2673, 16) & to_unsigned(6998, 16) & to_unsigned(31378, 16)),
    11 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(15181, 16) & to_unsigned(13645, 16) & to_unsigned(34501, 16) & to_unsigned(3393, 16) & to_unsigned(3840, 16) & to_unsigned(35227, 16) & to_unsigned(15562, 16) & to_unsigned(23615, 16) & to_unsigned(38342, 16) & to_unsigned(12139, 16) & to_unsigned(19471, 16) & to_unsigned(15483, 16)),
    12 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(13350, 16) & to_unsigned(6707, 16) & to_unsigned(23709, 16) & to_unsigned(37204, 16) & to_unsigned(25778, 16) & to_unsigned(21082, 16) & to_unsigned(7511, 16) & to_unsigned(14588, 16) & to_unsigned(10010, 16) & to_unsigned(21854, 16) & to_unsigned(28375, 16) & to_unsigned(33591, 16)),
    13 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(12514, 16) & to_unsigned(4695, 16) & to_unsigned(37190, 16) & to_unsigned(21379, 16) & to_unsigned(18723, 16) & to_unsigned(5802, 16) & to_unsigned(7182, 16) & to_unsigned(2529, 16) & to_unsigned(29936, 16) & to_unsigned(35860, 16) & to_unsigned(28338, 16) & to_unsigned(10835, 16)),
    14 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(34283, 16) & to_unsigned(25610, 16) & to_unsigned(33026, 16) & to_unsigned(31017, 16) & to_unsigned(21259, 16) & to_unsigned(2165, 16) & to_unsigned(21807, 16) & to_unsigned(37578, 16) & to_unsigned(1175, 16) & to_unsigned(16710, 16) & to_unsigned(21939, 16) & to_unsigned(30841, 16)),
    15 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(27292, 16) & to_unsigned(33730, 16) & to_unsigned(6836, 16) & to_unsigned(26476, 16) & to_unsigned(27539, 16) & to_unsigned(35784, 16) & to_unsigned(18245, 16) & to_unsigned(16394, 16) & to_unsigned(17939, 16) & to_unsigned(23094, 16) & to_unsigned(19216, 16) & to_unsigned(17432, 16)),
    16 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(11655, 16) & to_unsigned(6183, 16) & to_unsigned(38708, 16) & to_unsigned(28408, 16) & to_unsigned(35157, 16) & to_unsigned(17089, 16) & to_unsigned(13998, 16) & to_unsigned(36029, 16) & to_unsigned(15052, 16) & to_unsigned(16617, 16) & to_unsigned(5638, 16) & to_unsigned(36464, 16)),
    17 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(15693, 16) & to_unsigned(28923, 16) & to_unsigned(26245, 16) & to_unsigned(9432, 16) & to_unsigned(11675, 16) & to_unsigned(25720, 16) & to_unsigned(26405, 16) & to_unsigned(5838, 16) & to_unsigned(31851, 16) & to_unsigned(26898, 16) & to_unsigned(8090, 16) & to_unsigned(37037, 16)),
    18 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(24418, 16) & to_unsigned(27583, 16) & to_unsigned(7959, 16) & to_unsigned(35562, 16) & to_unsigned(37771, 16) & to_unsigned(17784, 16) & to_unsigned(11382, 16) & to_unsigned(11156, 16) & to_unsigned(37855, 16) & to_unsigned(7073, 16) & to_unsigned(21685, 16) & to_unsigned(34515, 16)),
    19 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(10977, 16) & to_unsigned(13633, 16) & to_unsigned(30969, 16) & to_unsigned(7516, 16) & to_unsigned(11943, 16) & to_unsigned(18199, 16) & to_unsigned(5231, 16) & to_unsigned(13825, 16) & to_unsigned(19589, 16) & to_unsigned(23661, 16) & to_unsigned(11150, 16) & to_unsigned(35602, 16)),
    20 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(19124, 16) & to_unsigned(30774, 16) & to_unsigned(6670, 16) & to_unsigned(37344, 16) & to_unsigned(16510, 16) & to_unsigned(26317, 16) & to_unsigned(23518, 16) & to_unsigned(22957, 16) & to_unsigned(6348, 16) & to_unsigned(34069, 16) & to_unsigned(8845, 16) & to_unsigned(20175, 16)),
    21 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(34985, 16) & to_unsigned(14441, 16) & to_unsigned(25668, 16) & to_unsigned(4116, 16) & to_unsigned(3019, 16) & to_unsigned(21049, 16) & to_unsigned(37308, 16) & to_unsigned(24551, 16) & to_unsigned(24727, 16) & to_unsigned(20104, 16) & to_unsigned(24850, 16) & to_unsigned(12114, 16)),
    22 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(38187, 16) & to_unsigned(28527, 16) & to_unsigned(13108, 16) & to_unsigned(13985, 16) & to_unsigned(1425, 16) & to_unsigned(21477, 16) & to_unsigned(30807, 16) & to_unsigned(8613, 16) & to_unsigned(26241, 16) & to_unsigned(33368, 16) & to_unsigned(35913, 16) & to_unsigned(32477, 16)),
    23 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(5903, 16) & to_unsigned(34390, 16) & to_unsigned(24641, 16) & to_unsigned(26556, 16) & to_unsigned(23007, 16) & to_unsigned(27305, 16) & to_unsigned(38247, 16) & to_unsigned(2621, 16) & to_unsigned(9122, 16) & to_unsigned(32806, 16) & to_unsigned(21554, 16) & to_unsigned(18685, 16)),
    24 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(17287, 16) & to_unsigned(27292, 16) & to_unsigned(19033, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    25 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(25796, 16) & to_unsigned(31795, 16) & to_unsigned(12152, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    26 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(12184, 16) & to_unsigned(35088, 16) & to_unsigned(31226, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    27 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(38263, 16) & to_unsigned(33386, 16) & to_unsigned(24892, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    28 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(23114, 16) & to_unsigned(37995, 16) & to_unsigned(29796, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    29 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(34336, 16) & to_unsigned(10551, 16) & to_unsigned(36245, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    30 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(35407, 16) & to_unsigned(175, 16) & to_unsigned(7203, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    31 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(14654, 16) & to_unsigned(38201, 16) & to_unsigned(22605, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    32 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(28404, 16) & to_unsigned(6595, 16) & to_unsigned(1018, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    33 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(19932, 16) & to_unsigned(3524, 16) & to_unsigned(29305, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    34 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(31749, 16) & to_unsigned(20247, 16) & to_unsigned(8128, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    35 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(18026, 16) & to_unsigned(36357, 16) & to_unsigned(26735, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    36 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7543, 16) & to_unsigned(29767, 16) & to_unsigned(13588, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    37 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(13333, 16) & to_unsigned(25965, 16) & to_unsigned(8463, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    38 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(14504, 16) & to_unsigned(36796, 16) & to_unsigned(19710, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    39 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4528, 16) & to_unsigned(25299, 16) & to_unsigned(7318, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    40 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(35091, 16) & to_unsigned(25550, 16) & to_unsigned(14798, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    41 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7824, 16) & to_unsigned(215, 16) & to_unsigned(1248, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    42 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(30848, 16) & to_unsigned(5362, 16) & to_unsigned(17291, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    43 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(28932, 16) & to_unsigned(30249, 16) & to_unsigned(27073, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    44 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(13062, 16) & to_unsigned(2103, 16) & to_unsigned(16206, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    45 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7129, 16) & to_unsigned(32062, 16) & to_unsigned(19612, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    46 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9512, 16) & to_unsigned(21936, 16) & to_unsigned(38833, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    47 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(35849, 16) & to_unsigned(33754, 16) & to_unsigned(23450, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    48 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(18705, 16) & to_unsigned(28656, 16) & to_unsigned(18111, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    49 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(22749, 16) & to_unsigned(27456, 16) & to_unsigned(32187, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    50 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(28229, 16) & to_unsigned(31684, 16) & to_unsigned(30160, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    51 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(15293, 16) & to_unsigned(8483, 16) & to_unsigned(28002, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    52 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(14880, 16) & to_unsigned(13334, 16) & to_unsigned(12584, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    53 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(28646, 16) & to_unsigned(2558, 16) & to_unsigned(19687, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    54 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6259, 16) & to_unsigned(4499, 16) & to_unsigned(26336, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    55 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(11952, 16) & to_unsigned(28386, 16) & to_unsigned(8405, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    56 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10609, 16) & to_unsigned(961, 16) & to_unsigned(7582, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    57 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10423, 16) & to_unsigned(13191, 16) & to_unsigned(26818, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    58 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(15922, 16) & to_unsigned(36654, 16) & to_unsigned(21450, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    59 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10492, 16) & to_unsigned(1532, 16) & to_unsigned(1205, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    60 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(30551, 16) & to_unsigned(36482, 16) & to_unsigned(22153, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    61 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5156, 16) & to_unsigned(11330, 16) & to_unsigned(34243, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    62 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(28616, 16) & to_unsigned(35369, 16) & to_unsigned(13322, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    63 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(8962, 16) & to_unsigned(1485, 16) & to_unsigned(21186, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    64 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(23541, 16) & to_unsigned(17445, 16) & to_unsigned(35561, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    65 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(33133, 16) & to_unsigned(11593, 16) & to_unsigned(19895, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    66 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(33917, 16) & to_unsigned(7863, 16) & to_unsigned(33651, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    67 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(20063, 16) & to_unsigned(28331, 16) & to_unsigned(10702, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    68 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(13195, 16) & to_unsigned(21107, 16) & to_unsigned(21859, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    69 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4364, 16) & to_unsigned(31137, 16) & to_unsigned(4804, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    70 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5585, 16) & to_unsigned(2037, 16) & to_unsigned(4830, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U')),
    71 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(30672, 16) & to_unsigned(16927, 16) & to_unsigned(14800, 16) & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U') & (15 downto 0 => 'U'))
  );

  -- From /home/souto/phase4ground/tables/ldpc/dvb/orig/dvb_64800_s2_b4_t2_a1.txt, table is 90x115 (1293.75 bytes)
  -- Resource estimation: 7 x 18 kB BRAMs or 4 x 36 kB BRAMs
  type dvb_64800_s2_b4_t2_a1_t is array (89 downto 0) of std_logic_vector(114 downto 0);

  constant DVB_64800_S2_B4_T2_A1_COLUMN_WIDTHS : integer_array_t := (0 => 3, 1 => 7, 2 => 15, 3 => 15, 4 => 15, 5 => 15, 6 => 15, 7 => 15, 8 => 15);

  constant DVB_64800_S2_B4_T2_A1 : dvb_64800_s2_b4_t2_a1_t := (
    0 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(54, 7) & to_unsigned(9318, 15) & to_unsigned(14392, 15) & to_unsigned(27561, 15) & to_unsigned(26909, 15) & to_unsigned(10219, 15) & to_unsigned(2534, 15) & to_unsigned(8597, 15)),
    1 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(55, 7) & to_unsigned(7263, 15) & to_unsigned(4635, 15) & to_unsigned(2530, 15) & to_unsigned(28130, 15) & to_unsigned(3033, 15) & to_unsigned(23830, 15) & to_unsigned(3651, 15)),
    2 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(56, 7) & to_unsigned(24731, 15) & to_unsigned(23583, 15) & to_unsigned(26036, 15) & to_unsigned(17299, 15) & to_unsigned(5750, 15) & to_unsigned(792, 15) & to_unsigned(9169, 15)),
    3 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(57, 7) & to_unsigned(5811, 15) & to_unsigned(26154, 15) & to_unsigned(18653, 15) & to_unsigned(11551, 15) & to_unsigned(15447, 15) & to_unsigned(13685, 15) & to_unsigned(16264, 15)),
    4 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(58, 7) & to_unsigned(12610, 15) & to_unsigned(11347, 15) & to_unsigned(28768, 15) & to_unsigned(2792, 15) & to_unsigned(3174, 15) & to_unsigned(29371, 15) & to_unsigned(12997, 15)),
    5 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(59, 7) & to_unsigned(16789, 15) & to_unsigned(16018, 15) & to_unsigned(21449, 15) & to_unsigned(6165, 15) & to_unsigned(21202, 15) & to_unsigned(15850, 15) & to_unsigned(3186, 15)),
    6 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(60, 7) & to_unsigned(31016, 15) & to_unsigned(21449, 15) & to_unsigned(17618, 15) & to_unsigned(6213, 15) & to_unsigned(12166, 15) & to_unsigned(8334, 15) & to_unsigned(18212, 15)),
    7 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(61, 7) & to_unsigned(22836, 15) & to_unsigned(14213, 15) & to_unsigned(11327, 15) & to_unsigned(5896, 15) & to_unsigned(718, 15) & to_unsigned(11727, 15) & to_unsigned(9308, 15)),
    8 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(62, 7) & to_unsigned(2091, 15) & to_unsigned(24941, 15) & to_unsigned(29966, 15) & to_unsigned(23634, 15) & to_unsigned(9013, 15) & to_unsigned(15587, 15) & to_unsigned(5444, 15)),
    9 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(63, 7) & to_unsigned(22207, 15) & to_unsigned(3983, 15) & to_unsigned(16904, 15) & to_unsigned(28534, 15) & to_unsigned(21415, 15) & to_unsigned(27524, 15) & to_unsigned(25912, 15)),
    10 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(64, 7) & to_unsigned(25687, 15) & to_unsigned(4501, 15) & to_unsigned(22193, 15) & to_unsigned(14665, 15) & to_unsigned(14798, 15) & to_unsigned(16158, 15) & to_unsigned(5491, 15)),
    11 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(65, 7) & to_unsigned(4520, 15) & to_unsigned(17094, 15) & to_unsigned(23397, 15) & to_unsigned(4264, 15) & to_unsigned(22370, 15) & to_unsigned(16941, 15) & to_unsigned(21526, 15)),
    12 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(66, 7) & to_unsigned(10490, 15) & to_unsigned(6182, 15) & to_unsigned(32370, 15) & to_unsigned(9597, 15) & to_unsigned(30841, 15) & to_unsigned(25954, 15) & to_unsigned(2762, 15)),
    13 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(67, 7) & to_unsigned(22120, 15) & to_unsigned(22865, 15) & to_unsigned(29870, 15) & to_unsigned(15147, 15) & to_unsigned(13668, 15) & to_unsigned(14955, 15) & to_unsigned(19235, 15)),
    14 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(68, 7) & to_unsigned(6689, 15) & to_unsigned(18408, 15) & to_unsigned(18346, 15) & to_unsigned(9918, 15) & to_unsigned(25746, 15) & to_unsigned(5443, 15) & to_unsigned(20645, 15)),
    15 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(69, 7) & to_unsigned(29982, 15) & to_unsigned(12529, 15) & to_unsigned(13858, 15) & to_unsigned(4746, 15) & to_unsigned(30370, 15) & to_unsigned(10023, 15) & to_unsigned(24828, 15)),
    16 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(70, 7) & to_unsigned(1262, 15) & to_unsigned(28032, 15) & to_unsigned(29888, 15) & to_unsigned(13063, 15) & to_unsigned(24033, 15) & to_unsigned(21951, 15) & to_unsigned(7863, 15)),
    17 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(71, 7) & to_unsigned(6594, 15) & to_unsigned(29642, 15) & to_unsigned(31451, 15) & to_unsigned(14831, 15) & to_unsigned(9509, 15) & to_unsigned(9335, 15) & to_unsigned(31552, 15)),
    18 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(72, 7) & to_unsigned(1358, 15) & to_unsigned(6454, 15) & to_unsigned(16633, 15) & to_unsigned(20354, 15) & to_unsigned(24598, 15) & to_unsigned(624, 15) & to_unsigned(5265, 15)),
    19 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(73, 7) & to_unsigned(19529, 15) & to_unsigned(295, 15) & to_unsigned(18011, 15) & to_unsigned(3080, 15) & to_unsigned(13364, 15) & to_unsigned(8032, 15) & to_unsigned(15323, 15)),
    20 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(74, 7) & to_unsigned(11981, 15) & to_unsigned(1510, 15) & to_unsigned(7960, 15) & to_unsigned(21462, 15) & to_unsigned(9129, 15) & to_unsigned(11370, 15) & to_unsigned(25741, 15)),
    21 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(75, 7) & to_unsigned(9276, 15) & to_unsigned(29656, 15) & to_unsigned(4543, 15) & to_unsigned(30699, 15) & to_unsigned(20646, 15) & to_unsigned(21921, 15) & to_unsigned(28050, 15)),
    22 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(76, 7) & to_unsigned(15975, 15) & to_unsigned(25634, 15) & to_unsigned(5520, 15) & to_unsigned(31119, 15) & to_unsigned(13715, 15) & to_unsigned(21949, 15) & to_unsigned(19605, 15)),
    23 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(77, 7) & to_unsigned(18688, 15) & to_unsigned(4608, 15) & to_unsigned(31755, 15) & to_unsigned(30165, 15) & to_unsigned(13103, 15) & to_unsigned(10706, 15) & to_unsigned(29224, 15)),
    24 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(78, 7) & to_unsigned(21514, 15) & to_unsigned(23117, 15) & to_unsigned(12245, 15) & to_unsigned(26035, 15) & to_unsigned(31656, 15) & to_unsigned(25631, 15) & to_unsigned(30699, 15)),
    25 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(79, 7) & to_unsigned(9674, 15) & to_unsigned(24966, 15) & to_unsigned(31285, 15) & to_unsigned(29908, 15) & to_unsigned(17042, 15) & to_unsigned(24588, 15) & to_unsigned(31857, 15)),
    26 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(80, 7) & to_unsigned(21856, 15) & to_unsigned(27777, 15) & to_unsigned(29919, 15) & to_unsigned(27000, 15) & to_unsigned(14897, 15) & to_unsigned(11409, 15) & to_unsigned(7122, 15)),
    27 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(81, 7) & to_unsigned(29773, 15) & to_unsigned(23310, 15) & to_unsigned(263, 15) & to_unsigned(4877, 15) & to_unsigned(28622, 15) & to_unsigned(20545, 15) & to_unsigned(22092, 15)),
    28 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(82, 7) & to_unsigned(15605, 15) & to_unsigned(5651, 15) & to_unsigned(21864, 15) & to_unsigned(3967, 15) & to_unsigned(14419, 15) & to_unsigned(22757, 15) & to_unsigned(15896, 15)),
    29 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(83, 7) & to_unsigned(30145, 15) & to_unsigned(1759, 15) & to_unsigned(10139, 15) & to_unsigned(29223, 15) & to_unsigned(26086, 15) & to_unsigned(10556, 15) & to_unsigned(5098, 15)),
    30 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(84, 7) & to_unsigned(18815, 15) & to_unsigned(16575, 15) & to_unsigned(2936, 15) & to_unsigned(24457, 15) & to_unsigned(26738, 15) & to_unsigned(6030, 15) & to_unsigned(505, 15)),
    31 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(85, 7) & to_unsigned(30326, 15) & to_unsigned(22298, 15) & to_unsigned(27562, 15) & to_unsigned(20131, 15) & to_unsigned(26390, 15) & to_unsigned(6247, 15) & to_unsigned(24791, 15)),
    32 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(86, 7) & to_unsigned(928, 15) & to_unsigned(29246, 15) & to_unsigned(21246, 15) & to_unsigned(12400, 15) & to_unsigned(15311, 15) & to_unsigned(32309, 15) & to_unsigned(18608, 15)),
    33 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(87, 7) & to_unsigned(20314, 15) & to_unsigned(6025, 15) & to_unsigned(26689, 15) & to_unsigned(16302, 15) & to_unsigned(2296, 15) & to_unsigned(3244, 15) & to_unsigned(19613, 15)),
    34 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(88, 7) & to_unsigned(6237, 15) & to_unsigned(11943, 15) & to_unsigned(22851, 15) & to_unsigned(15642, 15) & to_unsigned(23857, 15) & to_unsigned(15112, 15) & to_unsigned(20947, 15)),
    35 => std_logic_vector(to_unsigned(8, 3) & to_unsigned(89, 7) & to_unsigned(26403, 15) & to_unsigned(25168, 15) & to_unsigned(19038, 15) & to_unsigned(18384, 15) & to_unsigned(8882, 15) & to_unsigned(12719, 15) & to_unsigned(7093, 15)),
    36 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(0, 7) & to_unsigned(14567, 15) & to_unsigned(24965, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    37 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(1, 7) & to_unsigned(3908, 15) & to_unsigned(100, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    38 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(2, 7) & to_unsigned(10279, 15) & to_unsigned(240, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    39 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(3, 7) & to_unsigned(24102, 15) & to_unsigned(764, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    40 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(4, 7) & to_unsigned(12383, 15) & to_unsigned(4173, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    41 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(5, 7) & to_unsigned(13861, 15) & to_unsigned(15918, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    42 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(6, 7) & to_unsigned(21327, 15) & to_unsigned(1046, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    43 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(7, 7) & to_unsigned(5288, 15) & to_unsigned(14579, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    44 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(8, 7) & to_unsigned(28158, 15) & to_unsigned(8069, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    45 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(9, 7) & to_unsigned(16583, 15) & to_unsigned(11098, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    46 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(10, 7) & to_unsigned(16681, 15) & to_unsigned(28363, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    47 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(11, 7) & to_unsigned(13980, 15) & to_unsigned(24725, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    48 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(12, 7) & to_unsigned(32169, 15) & to_unsigned(17989, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    49 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(13, 7) & to_unsigned(10907, 15) & to_unsigned(2767, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    50 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(14, 7) & to_unsigned(21557, 15) & to_unsigned(3818, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    51 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(15, 7) & to_unsigned(26676, 15) & to_unsigned(12422, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    52 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(16, 7) & to_unsigned(7676, 15) & to_unsigned(8754, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    53 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(17, 7) & to_unsigned(14905, 15) & to_unsigned(20232, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    54 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(18, 7) & to_unsigned(15719, 15) & to_unsigned(24646, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    55 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(19, 7) & to_unsigned(31942, 15) & to_unsigned(8589, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    56 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(20, 7) & to_unsigned(19978, 15) & to_unsigned(27197, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    57 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(21, 7) & to_unsigned(27060, 15) & to_unsigned(15071, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    58 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(22, 7) & to_unsigned(6071, 15) & to_unsigned(26649, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    59 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(23, 7) & to_unsigned(10393, 15) & to_unsigned(11176, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    60 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(24, 7) & to_unsigned(9597, 15) & to_unsigned(13370, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    61 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(25, 7) & to_unsigned(7081, 15) & to_unsigned(17677, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    62 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(26, 7) & to_unsigned(1433, 15) & to_unsigned(19513, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    63 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(27, 7) & to_unsigned(26925, 15) & to_unsigned(9014, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    64 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(28, 7) & to_unsigned(19202, 15) & to_unsigned(8900, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    65 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(29, 7) & to_unsigned(18152, 15) & to_unsigned(30647, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    66 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(30, 7) & to_unsigned(20803, 15) & to_unsigned(1737, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    67 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(31, 7) & to_unsigned(11804, 15) & to_unsigned(25221, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    68 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(32, 7) & to_unsigned(31683, 15) & to_unsigned(17783, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    69 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(33, 7) & to_unsigned(29694, 15) & to_unsigned(9345, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    70 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(34, 7) & to_unsigned(12280, 15) & to_unsigned(26611, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    71 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(35, 7) & to_unsigned(6526, 15) & to_unsigned(26122, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    72 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(36, 7) & to_unsigned(26165, 15) & to_unsigned(11241, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    73 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(37, 7) & to_unsigned(7666, 15) & to_unsigned(26962, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    74 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(38, 7) & to_unsigned(16290, 15) & to_unsigned(8480, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    75 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(39, 7) & to_unsigned(11774, 15) & to_unsigned(10120, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    76 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(40, 7) & to_unsigned(30051, 15) & to_unsigned(30426, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    77 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(41, 7) & to_unsigned(1335, 15) & to_unsigned(15424, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    78 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(42, 7) & to_unsigned(6865, 15) & to_unsigned(17742, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    79 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(43, 7) & to_unsigned(31779, 15) & to_unsigned(12489, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    80 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(44, 7) & to_unsigned(32120, 15) & to_unsigned(21001, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    81 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(45, 7) & to_unsigned(14508, 15) & to_unsigned(6996, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    82 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(46, 7) & to_unsigned(979, 15) & to_unsigned(25024, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    83 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(47, 7) & to_unsigned(4554, 15) & to_unsigned(21896, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    84 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(48, 7) & to_unsigned(7989, 15) & to_unsigned(21777, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    85 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(49, 7) & to_unsigned(4972, 15) & to_unsigned(20661, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    86 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(50, 7) & to_unsigned(6612, 15) & to_unsigned(2730, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    87 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(51, 7) & to_unsigned(12742, 15) & to_unsigned(4418, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    88 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(52, 7) & to_unsigned(29194, 15) & to_unsigned(595, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    89 => std_logic_vector(to_unsigned(3, 3) & to_unsigned(53, 7) & to_unsigned(19267, 15) & to_unsigned(20113, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U'))
  );

  -- From /home/souto/phase4ground/tables/ldpc/dvb/orig/dvb_64800_s2_b5_t2_a2.txt, table is 108x184 (2484.0 bytes)
  -- Resource estimation: 11 x 18 kB BRAMs or 6 x 36 kB BRAMs
  type dvb_64800_s2_b5_t2_a2_t is array (107 downto 0) of std_logic_vector(183 downto 0);

  constant DVB_64800_S2_B5_T2_A2_COLUMN_WIDTHS : integer_array_t := (0 => 4, 1 => 15, 2 => 15, 3 => 15, 4 => 15, 5 => 15, 6 => 15, 7 => 15, 8 => 15, 9 => 15, 10 => 15, 11 => 15, 12 => 15);

  constant DVB_64800_S2_B5_T2_A2 : dvb_64800_s2_b5_t2_a2_t := (
    0 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(22422, 15) & to_unsigned(10282, 15) & to_unsigned(11626, 15) & to_unsigned(19997, 15) & to_unsigned(11161, 15) & to_unsigned(2922, 15) & to_unsigned(3122, 15) & to_unsigned(99, 15) & to_unsigned(5625, 15) & to_unsigned(17064, 15) & to_unsigned(8270, 15) & to_unsigned(179, 15)),
    1 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(25087, 15) & to_unsigned(16218, 15) & to_unsigned(17015, 15) & to_unsigned(828, 15) & to_unsigned(20041, 15) & to_unsigned(25656, 15) & to_unsigned(4186, 15) & to_unsigned(11629, 15) & to_unsigned(22599, 15) & to_unsigned(17305, 15) & to_unsigned(22515, 15) & to_unsigned(6463, 15)),
    2 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(11049, 15) & to_unsigned(22853, 15) & to_unsigned(25706, 15) & to_unsigned(14388, 15) & to_unsigned(5500, 15) & to_unsigned(19245, 15) & to_unsigned(8732, 15) & to_unsigned(2177, 15) & to_unsigned(13555, 15) & to_unsigned(11346, 15) & to_unsigned(17265, 15) & to_unsigned(3069, 15)),
    3 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(16581, 15) & to_unsigned(22225, 15) & to_unsigned(12563, 15) & to_unsigned(19717, 15) & to_unsigned(23577, 15) & to_unsigned(11555, 15) & to_unsigned(25496, 15) & to_unsigned(6853, 15) & to_unsigned(25403, 15) & to_unsigned(5218, 15) & to_unsigned(15925, 15) & to_unsigned(21766, 15)),
    4 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(16529, 15) & to_unsigned(14487, 15) & to_unsigned(7643, 15) & to_unsigned(10715, 15) & to_unsigned(17442, 15) & to_unsigned(11119, 15) & to_unsigned(5679, 15) & to_unsigned(14155, 15) & to_unsigned(24213, 15) & to_unsigned(21000, 15) & to_unsigned(1116, 15) & to_unsigned(15620, 15)),
    5 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(5340, 15) & to_unsigned(8636, 15) & to_unsigned(16693, 15) & to_unsigned(1434, 15) & to_unsigned(5635, 15) & to_unsigned(6516, 15) & to_unsigned(9482, 15) & to_unsigned(20189, 15) & to_unsigned(1066, 15) & to_unsigned(15013, 15) & to_unsigned(25361, 15) & to_unsigned(14243, 15)),
    6 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(18506, 15) & to_unsigned(22236, 15) & to_unsigned(20912, 15) & to_unsigned(8952, 15) & to_unsigned(5421, 15) & to_unsigned(15691, 15) & to_unsigned(6126, 15) & to_unsigned(21595, 15) & to_unsigned(500, 15) & to_unsigned(6904, 15) & to_unsigned(13059, 15) & to_unsigned(6802, 15)),
    7 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(8433, 15) & to_unsigned(4694, 15) & to_unsigned(5524, 15) & to_unsigned(14216, 15) & to_unsigned(3685, 15) & to_unsigned(19721, 15) & to_unsigned(25420, 15) & to_unsigned(9937, 15) & to_unsigned(23813, 15) & to_unsigned(9047, 15) & to_unsigned(25651, 15) & to_unsigned(16826, 15)),
    8 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(21500, 15) & to_unsigned(24814, 15) & to_unsigned(6344, 15) & to_unsigned(17382, 15) & to_unsigned(7064, 15) & to_unsigned(13929, 15) & to_unsigned(4004, 15) & to_unsigned(16552, 15) & to_unsigned(12818, 15) & to_unsigned(8720, 15) & to_unsigned(5286, 15) & to_unsigned(2206, 15)),
    9 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(22517, 15) & to_unsigned(2429, 15) & to_unsigned(19065, 15) & to_unsigned(2921, 15) & to_unsigned(21611, 15) & to_unsigned(1873, 15) & to_unsigned(7507, 15) & to_unsigned(5661, 15) & to_unsigned(23006, 15) & to_unsigned(23128, 15) & to_unsigned(20543, 15) & to_unsigned(19777, 15)),
    10 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(1770, 15) & to_unsigned(4636, 15) & to_unsigned(20900, 15) & to_unsigned(14931, 15) & to_unsigned(9247, 15) & to_unsigned(12340, 15) & to_unsigned(11008, 15) & to_unsigned(12966, 15) & to_unsigned(4471, 15) & to_unsigned(2731, 15) & to_unsigned(16445, 15) & to_unsigned(791, 15)),
    11 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(6635, 15) & to_unsigned(14556, 15) & to_unsigned(18865, 15) & to_unsigned(22421, 15) & to_unsigned(22124, 15) & to_unsigned(12697, 15) & to_unsigned(9803, 15) & to_unsigned(25485, 15) & to_unsigned(7744, 15) & to_unsigned(18254, 15) & to_unsigned(11313, 15) & to_unsigned(9004, 15)),
    12 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(19982, 15) & to_unsigned(23963, 15) & to_unsigned(18912, 15) & to_unsigned(7206, 15) & to_unsigned(12500, 15) & to_unsigned(4382, 15) & to_unsigned(20067, 15) & to_unsigned(6177, 15) & to_unsigned(21007, 15) & to_unsigned(1195, 15) & to_unsigned(23547, 15) & to_unsigned(24837, 15)),
    13 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(756, 15) & to_unsigned(11158, 15) & to_unsigned(14646, 15) & to_unsigned(20534, 15) & to_unsigned(3647, 15) & to_unsigned(17728, 15) & to_unsigned(11676, 15) & to_unsigned(11843, 15) & to_unsigned(12937, 15) & to_unsigned(4402, 15) & to_unsigned(8261, 15) & to_unsigned(22944, 15)),
    14 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(9306, 15) & to_unsigned(24009, 15) & to_unsigned(10012, 15) & to_unsigned(11081, 15) & to_unsigned(3746, 15) & to_unsigned(24325, 15) & to_unsigned(8060, 15) & to_unsigned(19826, 15) & to_unsigned(842, 15) & to_unsigned(8836, 15) & to_unsigned(2898, 15) & to_unsigned(5019, 15)),
    15 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(7575, 15) & to_unsigned(7455, 15) & to_unsigned(25244, 15) & to_unsigned(4736, 15) & to_unsigned(14400, 15) & to_unsigned(22981, 15) & to_unsigned(5543, 15) & to_unsigned(8006, 15) & to_unsigned(24203, 15) & to_unsigned(13053, 15) & to_unsigned(1120, 15) & to_unsigned(5128, 15)),
    16 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(3482, 15) & to_unsigned(9270, 15) & to_unsigned(13059, 15) & to_unsigned(15825, 15) & to_unsigned(7453, 15) & to_unsigned(23747, 15) & to_unsigned(3656, 15) & to_unsigned(24585, 15) & to_unsigned(16542, 15) & to_unsigned(17507, 15) & to_unsigned(22462, 15) & to_unsigned(14670, 15)),
    17 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(15627, 15) & to_unsigned(15290, 15) & to_unsigned(4198, 15) & to_unsigned(22748, 15) & to_unsigned(5842, 15) & to_unsigned(13395, 15) & to_unsigned(23918, 15) & to_unsigned(16985, 15) & to_unsigned(14929, 15) & to_unsigned(3726, 15) & to_unsigned(25350, 15) & to_unsigned(24157, 15)),
    18 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(24896, 15) & to_unsigned(16365, 15) & to_unsigned(16423, 15) & to_unsigned(13461, 15) & to_unsigned(16615, 15) & to_unsigned(8107, 15) & to_unsigned(24741, 15) & to_unsigned(3604, 15) & to_unsigned(25904, 15) & to_unsigned(8716, 15) & to_unsigned(9604, 15) & to_unsigned(20365, 15)),
    19 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(3729, 15) & to_unsigned(17245, 15) & to_unsigned(18448, 15) & to_unsigned(9862, 15) & to_unsigned(20831, 15) & to_unsigned(25326, 15) & to_unsigned(20517, 15) & to_unsigned(24618, 15) & to_unsigned(13282, 15) & to_unsigned(5099, 15) & to_unsigned(14183, 15) & to_unsigned(8804, 15)),
    20 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(16455, 15) & to_unsigned(17646, 15) & to_unsigned(15376, 15) & to_unsigned(18194, 15) & to_unsigned(25528, 15) & to_unsigned(1777, 15) & to_unsigned(6066, 15) & to_unsigned(21855, 15) & to_unsigned(14372, 15) & to_unsigned(12517, 15) & to_unsigned(4488, 15) & to_unsigned(17490, 15)),
    21 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(1400, 15) & to_unsigned(8135, 15) & to_unsigned(23375, 15) & to_unsigned(20879, 15) & to_unsigned(8476, 15) & to_unsigned(4084, 15) & to_unsigned(12936, 15) & to_unsigned(25536, 15) & to_unsigned(22309, 15) & to_unsigned(16582, 15) & to_unsigned(6402, 15) & to_unsigned(24360, 15)),
    22 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(25119, 15) & to_unsigned(23586, 15) & to_unsigned(128, 15) & to_unsigned(4761, 15) & to_unsigned(10443, 15) & to_unsigned(22536, 15) & to_unsigned(8607, 15) & to_unsigned(9752, 15) & to_unsigned(25446, 15) & to_unsigned(15053, 15) & to_unsigned(1856, 15) & to_unsigned(4040, 15)),
    23 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(377, 15) & to_unsigned(21160, 15) & to_unsigned(13474, 15) & to_unsigned(5451, 15) & to_unsigned(17170, 15) & to_unsigned(5938, 15) & to_unsigned(10256, 15) & to_unsigned(11972, 15) & to_unsigned(24210, 15) & to_unsigned(17833, 15) & to_unsigned(22047, 15) & to_unsigned(16108, 15)),
    24 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(13075, 15) & to_unsigned(9648, 15) & to_unsigned(24546, 15) & to_unsigned(13150, 15) & to_unsigned(23867, 15) & to_unsigned(7309, 15) & to_unsigned(19798, 15) & to_unsigned(2988, 15) & to_unsigned(16858, 15) & to_unsigned(4825, 15) & to_unsigned(23950, 15) & to_unsigned(15125, 15)),
    25 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(20526, 15) & to_unsigned(3553, 15) & to_unsigned(11525, 15) & to_unsigned(23366, 15) & to_unsigned(2452, 15) & to_unsigned(17626, 15) & to_unsigned(19265, 15) & to_unsigned(20172, 15) & to_unsigned(18060, 15) & to_unsigned(24593, 15) & to_unsigned(13255, 15) & to_unsigned(1552, 15)),
    26 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(18839, 15) & to_unsigned(21132, 15) & to_unsigned(20119, 15) & to_unsigned(15214, 15) & to_unsigned(14705, 15) & to_unsigned(7096, 15) & to_unsigned(10174, 15) & to_unsigned(5663, 15) & to_unsigned(18651, 15) & to_unsigned(19700, 15) & to_unsigned(12524, 15) & to_unsigned(14033, 15)),
    27 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(4127, 15) & to_unsigned(2971, 15) & to_unsigned(17499, 15) & to_unsigned(16287, 15) & to_unsigned(22368, 15) & to_unsigned(21463, 15) & to_unsigned(7943, 15) & to_unsigned(18880, 15) & to_unsigned(5567, 15) & to_unsigned(8047, 15) & to_unsigned(23363, 15) & to_unsigned(6797, 15)),
    28 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(10651, 15) & to_unsigned(24471, 15) & to_unsigned(14325, 15) & to_unsigned(4081, 15) & to_unsigned(7258, 15) & to_unsigned(4949, 15) & to_unsigned(7044, 15) & to_unsigned(1078, 15) & to_unsigned(797, 15) & to_unsigned(22910, 15) & to_unsigned(20474, 15) & to_unsigned(4318, 15)),
    29 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(21374, 15) & to_unsigned(13231, 15) & to_unsigned(22985, 15) & to_unsigned(5056, 15) & to_unsigned(3821, 15) & to_unsigned(23718, 15) & to_unsigned(14178, 15) & to_unsigned(9978, 15) & to_unsigned(19030, 15) & to_unsigned(23594, 15) & to_unsigned(8895, 15) & to_unsigned(25358, 15)),
    30 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(6199, 15) & to_unsigned(22056, 15) & to_unsigned(7749, 15) & to_unsigned(13310, 15) & to_unsigned(3999, 15) & to_unsigned(23697, 15) & to_unsigned(16445, 15) & to_unsigned(22636, 15) & to_unsigned(5225, 15) & to_unsigned(22437, 15) & to_unsigned(24153, 15) & to_unsigned(9442, 15)),
    31 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(7978, 15) & to_unsigned(12177, 15) & to_unsigned(2893, 15) & to_unsigned(20778, 15) & to_unsigned(3175, 15) & to_unsigned(8645, 15) & to_unsigned(11863, 15) & to_unsigned(24623, 15) & to_unsigned(10311, 15) & to_unsigned(25767, 15) & to_unsigned(17057, 15) & to_unsigned(3691, 15)),
    32 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(20473, 15) & to_unsigned(11294, 15) & to_unsigned(9914, 15) & to_unsigned(22815, 15) & to_unsigned(2574, 15) & to_unsigned(8439, 15) & to_unsigned(3699, 15) & to_unsigned(5431, 15) & to_unsigned(24840, 15) & to_unsigned(21908, 15) & to_unsigned(16088, 15) & to_unsigned(18244, 15)),
    33 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(8208, 15) & to_unsigned(5755, 15) & to_unsigned(19059, 15) & to_unsigned(8541, 15) & to_unsigned(24924, 15) & to_unsigned(6454, 15) & to_unsigned(11234, 15) & to_unsigned(10492, 15) & to_unsigned(16406, 15) & to_unsigned(10831, 15) & to_unsigned(11436, 15) & to_unsigned(9649, 15)),
    34 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(16264, 15) & to_unsigned(11275, 15) & to_unsigned(24953, 15) & to_unsigned(2347, 15) & to_unsigned(12667, 15) & to_unsigned(19190, 15) & to_unsigned(7257, 15) & to_unsigned(7174, 15) & to_unsigned(24819, 15) & to_unsigned(2938, 15) & to_unsigned(2522, 15) & to_unsigned(11749, 15)),
    35 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(3627, 15) & to_unsigned(5969, 15) & to_unsigned(13862, 15) & to_unsigned(1538, 15) & to_unsigned(23176, 15) & to_unsigned(6353, 15) & to_unsigned(2855, 15) & to_unsigned(17720, 15) & to_unsigned(2472, 15) & to_unsigned(7428, 15) & to_unsigned(573, 15) & to_unsigned(15036, 15)),
    36 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(0, 15) & to_unsigned(18539, 15) & to_unsigned(18661, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    37 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1, 15) & to_unsigned(10502, 15) & to_unsigned(3002, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    38 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(2, 15) & to_unsigned(9368, 15) & to_unsigned(10761, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    39 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3, 15) & to_unsigned(12299, 15) & to_unsigned(7828, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    40 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 15) & to_unsigned(15048, 15) & to_unsigned(13362, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    41 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 15) & to_unsigned(18444, 15) & to_unsigned(24640, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    42 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 15) & to_unsigned(20775, 15) & to_unsigned(19175, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    43 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 15) & to_unsigned(18970, 15) & to_unsigned(10971, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    44 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(8, 15) & to_unsigned(5329, 15) & to_unsigned(19982, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    45 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9, 15) & to_unsigned(11296, 15) & to_unsigned(18655, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    46 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10, 15) & to_unsigned(15046, 15) & to_unsigned(20659, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    47 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(11, 15) & to_unsigned(7300, 15) & to_unsigned(22140, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    48 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(12, 15) & to_unsigned(22029, 15) & to_unsigned(14477, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    49 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(13, 15) & to_unsigned(11129, 15) & to_unsigned(742, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    50 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(14, 15) & to_unsigned(13254, 15) & to_unsigned(13813, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    51 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(15, 15) & to_unsigned(19234, 15) & to_unsigned(13273, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    52 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(16, 15) & to_unsigned(6079, 15) & to_unsigned(21122, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    53 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(17, 15) & to_unsigned(22782, 15) & to_unsigned(5828, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    54 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(18, 15) & to_unsigned(19775, 15) & to_unsigned(4247, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    55 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(19, 15) & to_unsigned(1660, 15) & to_unsigned(19413, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    56 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(20, 15) & to_unsigned(4403, 15) & to_unsigned(3649, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    57 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(21, 15) & to_unsigned(13371, 15) & to_unsigned(25851, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    58 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(22, 15) & to_unsigned(22770, 15) & to_unsigned(21784, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    59 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(23, 15) & to_unsigned(10757, 15) & to_unsigned(14131, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    60 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(24, 15) & to_unsigned(16071, 15) & to_unsigned(21617, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    61 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(25, 15) & to_unsigned(6393, 15) & to_unsigned(3725, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    62 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(26, 15) & to_unsigned(597, 15) & to_unsigned(19968, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    63 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(27, 15) & to_unsigned(5743, 15) & to_unsigned(8084, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    64 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(28, 15) & to_unsigned(6770, 15) & to_unsigned(9548, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    65 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(29, 15) & to_unsigned(4285, 15) & to_unsigned(17542, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    66 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(30, 15) & to_unsigned(13568, 15) & to_unsigned(22599, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    67 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(31, 15) & to_unsigned(1786, 15) & to_unsigned(4617, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    68 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(32, 15) & to_unsigned(23238, 15) & to_unsigned(11648, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    69 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(33, 15) & to_unsigned(19627, 15) & to_unsigned(2030, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    70 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(34, 15) & to_unsigned(13601, 15) & to_unsigned(13458, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    71 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(35, 15) & to_unsigned(13740, 15) & to_unsigned(17328, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    72 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(36, 15) & to_unsigned(25012, 15) & to_unsigned(13944, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    73 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(37, 15) & to_unsigned(22513, 15) & to_unsigned(6687, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    74 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(38, 15) & to_unsigned(4934, 15) & to_unsigned(12587, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    75 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(39, 15) & to_unsigned(21197, 15) & to_unsigned(5133, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    76 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(40, 15) & to_unsigned(22705, 15) & to_unsigned(6938, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    77 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(41, 15) & to_unsigned(7534, 15) & to_unsigned(24633, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    78 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(42, 15) & to_unsigned(24400, 15) & to_unsigned(12797, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    79 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(43, 15) & to_unsigned(21911, 15) & to_unsigned(25712, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    80 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(44, 15) & to_unsigned(12039, 15) & to_unsigned(1140, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    81 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(45, 15) & to_unsigned(24306, 15) & to_unsigned(1021, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    82 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(46, 15) & to_unsigned(14012, 15) & to_unsigned(20747, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    83 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(47, 15) & to_unsigned(11265, 15) & to_unsigned(15219, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    84 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(48, 15) & to_unsigned(4670, 15) & to_unsigned(15531, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    85 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(49, 15) & to_unsigned(9417, 15) & to_unsigned(14359, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    86 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(50, 15) & to_unsigned(2415, 15) & to_unsigned(6504, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    87 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(51, 15) & to_unsigned(24964, 15) & to_unsigned(24690, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    88 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(52, 15) & to_unsigned(14443, 15) & to_unsigned(8816, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    89 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(53, 15) & to_unsigned(6926, 15) & to_unsigned(1291, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    90 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(54, 15) & to_unsigned(6209, 15) & to_unsigned(20806, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    91 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(55, 15) & to_unsigned(13915, 15) & to_unsigned(4079, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    92 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(56, 15) & to_unsigned(24410, 15) & to_unsigned(13196, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    93 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(57, 15) & to_unsigned(13505, 15) & to_unsigned(6117, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    94 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(58, 15) & to_unsigned(9869, 15) & to_unsigned(8220, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    95 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(59, 15) & to_unsigned(1570, 15) & to_unsigned(6044, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    96 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(60, 15) & to_unsigned(25780, 15) & to_unsigned(17387, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    97 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(61, 15) & to_unsigned(20671, 15) & to_unsigned(24913, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    98 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(62, 15) & to_unsigned(24558, 15) & to_unsigned(20591, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    99 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(63, 15) & to_unsigned(12402, 15) & to_unsigned(3702, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    100 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(64, 15) & to_unsigned(8314, 15) & to_unsigned(1357, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    101 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(65, 15) & to_unsigned(20071, 15) & to_unsigned(14616, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    102 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(66, 15) & to_unsigned(17014, 15) & to_unsigned(3688, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    103 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(67, 15) & to_unsigned(19837, 15) & to_unsigned(946, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    104 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(68, 15) & to_unsigned(15195, 15) & to_unsigned(12136, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    105 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(69, 15) & to_unsigned(7758, 15) & to_unsigned(22808, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    106 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(70, 15) & to_unsigned(3564, 15) & to_unsigned(2925, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    107 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(71, 15) & to_unsigned(3434, 15) & to_unsigned(7769, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U'))
  );

  -- From /home/souto/phase4ground/tables/ldpc/dvb/orig/dvb_64800_s2_b6.txt, table is 120x189 (2835.0 bytes)
  -- Resource estimation: 11 x 18 kB BRAMs or 6 x 36 kB BRAMs
  type dvb_64800_s2_b6_t is array (119 downto 0) of std_logic_vector(188 downto 0);

  constant DVB_64800_S2_B6_COLUMN_WIDTHS : integer_array_t := (0 => 4, 1 => 6, 2 => 15, 3 => 15, 4 => 15, 5 => 15, 6 => 15, 7 => 15, 8 => 14, 9 => 15, 10 => 15, 11 => 15, 12 => 15, 13 => 15);

  constant DVB_64800_S2_B6 : dvb_64800_s2_b6_t := (
    0 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(0, 6) & to_unsigned(10491, 15) & to_unsigned(16043, 15) & to_unsigned(506, 15) & to_unsigned(12826, 15) & to_unsigned(8065, 15) & to_unsigned(8226, 15) & to_unsigned(2767, 14) & to_unsigned(240, 15) & to_unsigned(18673, 15) & to_unsigned(9279, 15) & to_unsigned(10579, 15) & to_unsigned(20928, 15)),
    1 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(1, 6) & to_unsigned(17819, 15) & to_unsigned(8313, 15) & to_unsigned(6433, 15) & to_unsigned(6224, 15) & to_unsigned(5120, 15) & to_unsigned(5824, 15) & to_unsigned(12812, 14) & to_unsigned(17187, 15) & to_unsigned(9940, 15) & to_unsigned(13447, 15) & to_unsigned(13825, 15) & to_unsigned(18483, 15)),
    2 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(2, 6) & to_unsigned(17957, 15) & to_unsigned(6024, 15) & to_unsigned(8681, 15) & to_unsigned(18628, 15) & to_unsigned(12794, 15) & to_unsigned(5915, 15) & to_unsigned(14576, 14) & to_unsigned(10970, 15) & to_unsigned(12064, 15) & to_unsigned(20437, 15) & to_unsigned(4455, 15) & to_unsigned(7151, 15)),
    3 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(3, 6) & to_unsigned(19777, 15) & to_unsigned(6183, 15) & to_unsigned(9972, 15) & to_unsigned(14536, 15) & to_unsigned(8182, 15) & to_unsigned(17749, 15) & to_unsigned(11341, 14) & to_unsigned(5556, 15) & to_unsigned(4379, 15) & to_unsigned(17434, 15) & to_unsigned(15477, 15) & to_unsigned(18532, 15)),
    4 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(4, 6) & to_unsigned(4651, 15) & to_unsigned(19689, 15) & to_unsigned(1608, 15) & to_unsigned(659, 15) & to_unsigned(16707, 15) & to_unsigned(14335, 15) & to_unsigned(6143, 14) & to_unsigned(3058, 15) & to_unsigned(14618, 15) & to_unsigned(17894, 15) & to_unsigned(20684, 15) & to_unsigned(5306, 15)),
    5 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(5, 6) & to_unsigned(9778, 15) & to_unsigned(2552, 15) & to_unsigned(12096, 15) & to_unsigned(12369, 15) & to_unsigned(15198, 15) & to_unsigned(16890, 15) & to_unsigned(4851, 14) & to_unsigned(3109, 15) & to_unsigned(1700, 15) & to_unsigned(18725, 15) & to_unsigned(1997, 15) & to_unsigned(15882, 15)),
    6 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(6, 6) & to_unsigned(486, 15) & to_unsigned(6111, 15) & to_unsigned(13743, 15) & to_unsigned(11537, 15) & to_unsigned(5591, 15) & to_unsigned(7433, 15) & to_unsigned(15227, 14) & to_unsigned(14145, 15) & to_unsigned(1483, 15) & to_unsigned(3887, 15) & to_unsigned(17431, 15) & to_unsigned(12430, 15)),
    7 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(7, 6) & to_unsigned(20647, 15) & to_unsigned(14311, 15) & to_unsigned(11734, 15) & to_unsigned(4180, 15) & to_unsigned(8110, 15) & to_unsigned(5525, 15) & to_unsigned(12141, 14) & to_unsigned(15761, 15) & to_unsigned(18661, 15) & to_unsigned(18441, 15) & to_unsigned(10569, 15) & to_unsigned(8192, 15)),
    8 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(8, 6) & to_unsigned(3791, 15) & to_unsigned(14759, 15) & to_unsigned(15264, 15) & to_unsigned(19918, 15) & to_unsigned(10132, 15) & to_unsigned(9062, 15) & to_unsigned(10010, 14) & to_unsigned(12786, 15) & to_unsigned(10675, 15) & to_unsigned(9682, 15) & to_unsigned(19246, 15) & to_unsigned(5454, 15)),
    9 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(9, 6) & to_unsigned(19525, 15) & to_unsigned(9485, 15) & to_unsigned(7777, 15) & to_unsigned(19999, 15) & to_unsigned(8378, 15) & to_unsigned(9209, 15) & to_unsigned(3163, 14) & to_unsigned(20232, 15) & to_unsigned(6690, 15) & to_unsigned(16518, 15) & to_unsigned(716, 15) & to_unsigned(7353, 15)),
    10 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(10, 6) & to_unsigned(4588, 15) & to_unsigned(6709, 15) & to_unsigned(20202, 15) & to_unsigned(10905, 15) & to_unsigned(915, 15) & to_unsigned(4317, 15) & to_unsigned(11073, 14) & to_unsigned(13576, 15) & to_unsigned(16433, 15) & to_unsigned(368, 15) & to_unsigned(3508, 15) & to_unsigned(21171, 15)),
    11 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(11, 6) & to_unsigned(14072, 15) & to_unsigned(4033, 15) & to_unsigned(19959, 15) & to_unsigned(12608, 15) & to_unsigned(631, 15) & to_unsigned(19494, 15) & to_unsigned(14160, 14) & to_unsigned(8249, 15) & to_unsigned(10223, 15) & to_unsigned(21504, 15) & to_unsigned(12395, 15) & to_unsigned(4322, 15)),
    12 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(12, 6) & to_unsigned(13800, 15) & to_unsigned(14161, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    13 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(13, 6) & to_unsigned(2948, 15) & to_unsigned(9647, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    14 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(14, 6) & to_unsigned(14693, 15) & to_unsigned(16027, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    15 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(15, 6) & to_unsigned(20506, 15) & to_unsigned(11082, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    16 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(16, 6) & to_unsigned(1143, 15) & to_unsigned(9020, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    17 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(17, 6) & to_unsigned(13501, 15) & to_unsigned(4014, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    18 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(18, 6) & to_unsigned(1548, 15) & to_unsigned(2190, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    19 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(19, 6) & to_unsigned(12216, 15) & to_unsigned(21556, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    20 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(20, 6) & to_unsigned(2095, 15) & to_unsigned(19897, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    21 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(21, 6) & to_unsigned(4189, 15) & to_unsigned(7958, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    22 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(22, 6) & to_unsigned(15940, 15) & to_unsigned(10048, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    23 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(23, 6) & to_unsigned(515, 15) & to_unsigned(12614, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    24 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(24, 6) & to_unsigned(8501, 15) & to_unsigned(8450, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    25 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(25, 6) & to_unsigned(17595, 15) & to_unsigned(16784, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    26 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(26, 6) & to_unsigned(5913, 15) & to_unsigned(8495, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    27 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(27, 6) & to_unsigned(16394, 15) & to_unsigned(10423, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    28 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(28, 6) & to_unsigned(7409, 15) & to_unsigned(6981, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    29 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(29, 6) & to_unsigned(6678, 15) & to_unsigned(15939, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    30 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(30, 6) & to_unsigned(20344, 15) & to_unsigned(12987, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    31 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(31, 6) & to_unsigned(2510, 15) & to_unsigned(14588, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    32 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(32, 6) & to_unsigned(17918, 15) & to_unsigned(6655, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    33 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(33, 6) & to_unsigned(6703, 15) & to_unsigned(19451, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    34 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(34, 6) & to_unsigned(496, 15) & to_unsigned(4217, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    35 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(35, 6) & to_unsigned(7290, 15) & to_unsigned(5766, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    36 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(36, 6) & to_unsigned(10521, 15) & to_unsigned(8925, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    37 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(37, 6) & to_unsigned(20379, 15) & to_unsigned(11905, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    38 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(38, 6) & to_unsigned(4090, 15) & to_unsigned(5838, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    39 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(39, 6) & to_unsigned(19082, 15) & to_unsigned(17040, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    40 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(40, 6) & to_unsigned(20233, 15) & to_unsigned(12352, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    41 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(41, 6) & to_unsigned(19365, 15) & to_unsigned(19546, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    42 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(42, 6) & to_unsigned(6249, 15) & to_unsigned(19030, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    43 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(43, 6) & to_unsigned(11037, 15) & to_unsigned(19193, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    44 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(44, 6) & to_unsigned(19760, 15) & to_unsigned(11772, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    45 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(45, 6) & to_unsigned(19644, 15) & to_unsigned(7428, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    46 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(46, 6) & to_unsigned(16076, 15) & to_unsigned(3521, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    47 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(47, 6) & to_unsigned(11779, 15) & to_unsigned(21062, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    48 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(48, 6) & to_unsigned(13062, 15) & to_unsigned(9682, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    49 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(49, 6) & to_unsigned(8934, 15) & to_unsigned(5217, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    50 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(50, 6) & to_unsigned(11087, 15) & to_unsigned(3319, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    51 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(51, 6) & to_unsigned(18892, 15) & to_unsigned(4356, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    52 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(52, 6) & to_unsigned(7894, 15) & to_unsigned(3898, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    53 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(53, 6) & to_unsigned(5963, 15) & to_unsigned(4360, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    54 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(54, 6) & to_unsigned(7346, 15) & to_unsigned(11726, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    55 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(55, 6) & to_unsigned(5182, 15) & to_unsigned(5609, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    56 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(56, 6) & to_unsigned(2412, 15) & to_unsigned(17295, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    57 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(57, 6) & to_unsigned(9845, 15) & to_unsigned(20494, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    58 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(58, 6) & to_unsigned(6687, 15) & to_unsigned(1864, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    59 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(59, 6) & to_unsigned(20564, 15) & to_unsigned(5216, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    60 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(0, 6) & to_unsigned(18226, 15) & to_unsigned(17207, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    61 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1, 6) & to_unsigned(9380, 15) & to_unsigned(8266, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    62 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(2, 6) & to_unsigned(7073, 15) & to_unsigned(3065, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    63 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3, 6) & to_unsigned(18252, 15) & to_unsigned(13437, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    64 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 6) & to_unsigned(9161, 15) & to_unsigned(15642, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    65 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 6) & to_unsigned(10714, 15) & to_unsigned(10153, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    66 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 6) & to_unsigned(11585, 15) & to_unsigned(9078, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    67 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 6) & to_unsigned(5359, 15) & to_unsigned(9418, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    68 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(8, 6) & to_unsigned(9024, 15) & to_unsigned(9515, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    69 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9, 6) & to_unsigned(1206, 15) & to_unsigned(16354, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    70 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10, 6) & to_unsigned(14994, 15) & to_unsigned(1102, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    71 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(11, 6) & to_unsigned(9375, 15) & to_unsigned(20796, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    72 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(12, 6) & to_unsigned(15964, 15) & to_unsigned(6027, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    73 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(13, 6) & to_unsigned(14789, 15) & to_unsigned(6452, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    74 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(14, 6) & to_unsigned(8002, 15) & to_unsigned(18591, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    75 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(15, 6) & to_unsigned(14742, 15) & to_unsigned(14089, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    76 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(16, 6) & to_unsigned(253, 15) & to_unsigned(3045, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    77 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(17, 6) & to_unsigned(1274, 15) & to_unsigned(19286, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    78 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(18, 6) & to_unsigned(14777, 15) & to_unsigned(2044, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    79 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(19, 6) & to_unsigned(13920, 15) & to_unsigned(9900, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    80 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(20, 6) & to_unsigned(452, 15) & to_unsigned(7374, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    81 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(21, 6) & to_unsigned(18206, 15) & to_unsigned(9921, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    82 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(22, 6) & to_unsigned(6131, 15) & to_unsigned(5414, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    83 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(23, 6) & to_unsigned(10077, 15) & to_unsigned(9726, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    84 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(24, 6) & to_unsigned(12045, 15) & to_unsigned(5479, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    85 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(25, 6) & to_unsigned(4322, 15) & to_unsigned(7990, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    86 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(26, 6) & to_unsigned(15616, 15) & to_unsigned(5550, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    87 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(27, 6) & to_unsigned(15561, 15) & to_unsigned(10661, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    88 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(28, 6) & to_unsigned(20718, 15) & to_unsigned(7387, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    89 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(29, 6) & to_unsigned(2518, 15) & to_unsigned(18804, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    90 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(30, 6) & to_unsigned(8984, 15) & to_unsigned(2600, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    91 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(31, 6) & to_unsigned(6516, 15) & to_unsigned(17909, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    92 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(32, 6) & to_unsigned(11148, 15) & to_unsigned(98, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    93 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(33, 6) & to_unsigned(20559, 15) & to_unsigned(3704, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    94 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(34, 6) & to_unsigned(7510, 15) & to_unsigned(1569, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    95 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(35, 6) & to_unsigned(16000, 15) & to_unsigned(11692, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    96 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(36, 6) & to_unsigned(9147, 15) & to_unsigned(10303, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    97 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(37, 6) & to_unsigned(16650, 15) & to_unsigned(191, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    98 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(38, 6) & to_unsigned(15577, 15) & to_unsigned(18685, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    99 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(39, 6) & to_unsigned(17167, 15) & to_unsigned(20917, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    100 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(40, 6) & to_unsigned(4256, 15) & to_unsigned(3391, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    101 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(41, 6) & to_unsigned(20092, 15) & to_unsigned(17219, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    102 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(42, 6) & to_unsigned(9218, 15) & to_unsigned(5056, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    103 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(43, 6) & to_unsigned(18429, 15) & to_unsigned(8472, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    104 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(44, 6) & to_unsigned(12093, 15) & to_unsigned(20753, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    105 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(45, 6) & to_unsigned(16345, 15) & to_unsigned(12748, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    106 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(46, 6) & to_unsigned(16023, 15) & to_unsigned(11095, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    107 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(47, 6) & to_unsigned(5048, 15) & to_unsigned(17595, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    108 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(48, 6) & to_unsigned(18995, 15) & to_unsigned(4817, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    109 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(49, 6) & to_unsigned(16483, 15) & to_unsigned(3536, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    110 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(50, 6) & to_unsigned(1439, 15) & to_unsigned(16148, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    111 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(51, 6) & to_unsigned(3661, 15) & to_unsigned(3039, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    112 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(52, 6) & to_unsigned(19010, 15) & to_unsigned(18121, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    113 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(53, 6) & to_unsigned(8968, 15) & to_unsigned(11793, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    114 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(54, 6) & to_unsigned(13427, 15) & to_unsigned(18003, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    115 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(55, 6) & to_unsigned(5303, 15) & to_unsigned(3083, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    116 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(56, 6) & to_unsigned(531, 15) & to_unsigned(16668, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    117 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(57, 6) & to_unsigned(4771, 15) & to_unsigned(6722, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    118 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(58, 6) & to_unsigned(5695, 15) & to_unsigned(7960, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U')),
    119 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(59, 6) & to_unsigned(3589, 15) & to_unsigned(14630, 15) & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (13 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U') & (14 downto 0 => 'U'))
  );

  -- From /home/souto/phase4ground/tables/ldpc/dvb/orig/dvb_64800_s2_b7_t2_a4.txt, table is 135x164 (2767.5 bytes)
  -- Resource estimation: 10 x 18 kB BRAMs or 5 x 36 kB BRAMs
  type dvb_64800_s2_b7_t2_a4_t is array (134 downto 0) of std_logic_vector(163 downto 0);

  constant DVB_64800_S2_B7_T2_A4_COLUMN_WIDTHS : integer_array_t := (0 => 4, 1 => 6, 2 => 14, 3 => 14, 4 => 14, 5 => 14, 6 => 14, 7 => 14, 8 => 14, 9 => 14, 10 => 14, 11 => 14, 12 => 14);

  constant DVB_64800_S2_B7_T2_A4 : dvb_64800_s2_b7_t2_a4_t := (
    0 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(0, 6) & to_unsigned(6385, 14) & to_unsigned(7901, 14) & to_unsigned(14611, 14) & to_unsigned(13389, 14) & to_unsigned(11200, 14) & to_unsigned(3252, 14) & to_unsigned(5243, 14) & to_unsigned(2504, 14) & to_unsigned(2722, 14) & to_unsigned(821, 14) & to_unsigned(7374, 14)),
    1 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(1, 6) & to_unsigned(11359, 14) & to_unsigned(2698, 14) & to_unsigned(357, 14) & to_unsigned(13824, 14) & to_unsigned(12772, 14) & to_unsigned(7244, 14) & to_unsigned(6752, 14) & to_unsigned(15310, 14) & to_unsigned(852, 14) & to_unsigned(2001, 14) & to_unsigned(11417, 14)),
    2 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(2, 6) & to_unsigned(7862, 14) & to_unsigned(7977, 14) & to_unsigned(6321, 14) & to_unsigned(13612, 14) & to_unsigned(12197, 14) & to_unsigned(14449, 14) & to_unsigned(15137, 14) & to_unsigned(13860, 14) & to_unsigned(1708, 14) & to_unsigned(6399, 14) & to_unsigned(13444, 14)),
    3 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(3, 6) & to_unsigned(1560, 14) & to_unsigned(11804, 14) & to_unsigned(6975, 14) & to_unsigned(13292, 14) & to_unsigned(3646, 14) & to_unsigned(3812, 14) & to_unsigned(8772, 14) & to_unsigned(7306, 14) & to_unsigned(5795, 14) & to_unsigned(14327, 14) & to_unsigned(7866, 14)),
    4 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(4, 6) & to_unsigned(7626, 14) & to_unsigned(11407, 14) & to_unsigned(14599, 14) & to_unsigned(9689, 14) & to_unsigned(1628, 14) & to_unsigned(2113, 14) & to_unsigned(10809, 14) & to_unsigned(9283, 14) & to_unsigned(1230, 14) & to_unsigned(15241, 14) & to_unsigned(4870, 14)),
    5 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(5, 6) & to_unsigned(1610, 14) & to_unsigned(5699, 14) & to_unsigned(15876, 14) & to_unsigned(9446, 14) & to_unsigned(12515, 14) & to_unsigned(1400, 14) & to_unsigned(6303, 14) & to_unsigned(5411, 14) & to_unsigned(14181, 14) & to_unsigned(13925, 14) & to_unsigned(7358, 14)),
    6 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(6, 6) & to_unsigned(4059, 14) & to_unsigned(8836, 14) & to_unsigned(3405, 14) & to_unsigned(7853, 14) & to_unsigned(7992, 14) & to_unsigned(15336, 14) & to_unsigned(5970, 14) & to_unsigned(10368, 14) & to_unsigned(10278, 14) & to_unsigned(9675, 14) & to_unsigned(4651, 14)),
    7 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(7, 6) & to_unsigned(4441, 14) & to_unsigned(3963, 14) & to_unsigned(9153, 14) & to_unsigned(2109, 14) & to_unsigned(12683, 14) & to_unsigned(7459, 14) & to_unsigned(12030, 14) & to_unsigned(12221, 14) & to_unsigned(629, 14) & to_unsigned(15212, 14) & to_unsigned(406, 14)),
    8 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(8, 6) & to_unsigned(6007, 14) & to_unsigned(8411, 14) & to_unsigned(5771, 14) & to_unsigned(3497, 14) & to_unsigned(543, 14) & to_unsigned(14202, 14) & to_unsigned(875, 14) & to_unsigned(9186, 14) & to_unsigned(6235, 14) & to_unsigned(13908, 14) & to_unsigned(3563, 14)),
    9 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(9, 6) & to_unsigned(3232, 14) & to_unsigned(6625, 14) & to_unsigned(4795, 14) & to_unsigned(546, 14) & to_unsigned(9781, 14) & to_unsigned(2071, 14) & to_unsigned(7312, 14) & to_unsigned(3399, 14) & to_unsigned(7250, 14) & to_unsigned(4932, 14) & to_unsigned(12652, 14)),
    10 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(10, 6) & to_unsigned(8820, 14) & to_unsigned(10088, 14) & to_unsigned(11090, 14) & to_unsigned(7069, 14) & to_unsigned(6585, 14) & to_unsigned(13134, 14) & to_unsigned(10158, 14) & to_unsigned(7183, 14) & to_unsigned(488, 14) & to_unsigned(7455, 14) & to_unsigned(9238, 14)),
    11 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(11, 6) & to_unsigned(1903, 14) & to_unsigned(10818, 14) & to_unsigned(119, 14) & to_unsigned(215, 14) & to_unsigned(7558, 14) & to_unsigned(11046, 14) & to_unsigned(10615, 14) & to_unsigned(11545, 14) & to_unsigned(14784, 14) & to_unsigned(7961, 14) & to_unsigned(15619, 14)),
    12 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(12, 6) & to_unsigned(3655, 14) & to_unsigned(8736, 14) & to_unsigned(4917, 14) & to_unsigned(15874, 14) & to_unsigned(5129, 14) & to_unsigned(2134, 14) & to_unsigned(15944, 14) & to_unsigned(14768, 14) & to_unsigned(7150, 14) & to_unsigned(2692, 14) & to_unsigned(1469, 14)),
    13 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(13, 6) & to_unsigned(8316, 14) & to_unsigned(3820, 14) & to_unsigned(505, 14) & to_unsigned(8923, 14) & to_unsigned(6757, 14) & to_unsigned(806, 14) & to_unsigned(7957, 14) & to_unsigned(4216, 14) & to_unsigned(15589, 14) & to_unsigned(13244, 14) & to_unsigned(2622, 14)),
    14 => std_logic_vector(to_unsigned(12, 4) & to_unsigned(14, 6) & to_unsigned(14463, 14) & to_unsigned(4852, 14) & to_unsigned(15733, 14) & to_unsigned(3041, 14) & to_unsigned(11193, 14) & to_unsigned(12860, 14) & to_unsigned(13673, 14) & to_unsigned(8152, 14) & to_unsigned(6551, 14) & to_unsigned(15108, 14) & to_unsigned(8758, 14)),
    15 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(15, 6) & to_unsigned(3149, 14) & to_unsigned(11981, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    16 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(16, 6) & to_unsigned(13416, 14) & to_unsigned(6906, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    17 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(17, 6) & to_unsigned(13098, 14) & to_unsigned(13352, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    18 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(18, 6) & to_unsigned(2009, 14) & to_unsigned(14460, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    19 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(19, 6) & to_unsigned(7207, 14) & to_unsigned(4314, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    20 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(20, 6) & to_unsigned(3312, 14) & to_unsigned(3945, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    21 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(21, 6) & to_unsigned(4418, 14) & to_unsigned(6248, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    22 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(22, 6) & to_unsigned(2669, 14) & to_unsigned(13975, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    23 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(23, 6) & to_unsigned(7571, 14) & to_unsigned(9023, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    24 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(24, 6) & to_unsigned(14172, 14) & to_unsigned(2967, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    25 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(25, 6) & to_unsigned(7271, 14) & to_unsigned(7138, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    26 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(26, 6) & to_unsigned(6135, 14) & to_unsigned(13670, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    27 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(27, 6) & to_unsigned(7490, 14) & to_unsigned(14559, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    28 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(28, 6) & to_unsigned(8657, 14) & to_unsigned(2466, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    29 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(29, 6) & to_unsigned(8599, 14) & to_unsigned(12834, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    30 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(30, 6) & to_unsigned(3470, 14) & to_unsigned(3152, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    31 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(31, 6) & to_unsigned(13917, 14) & to_unsigned(4365, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    32 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(32, 6) & to_unsigned(6024, 14) & to_unsigned(13730, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    33 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(33, 6) & to_unsigned(10973, 14) & to_unsigned(14182, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    34 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(34, 6) & to_unsigned(2464, 14) & to_unsigned(13167, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    35 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(35, 6) & to_unsigned(5281, 14) & to_unsigned(15049, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    36 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(36, 6) & to_unsigned(1103, 14) & to_unsigned(1849, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    37 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(37, 6) & to_unsigned(2058, 14) & to_unsigned(1069, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    38 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(38, 6) & to_unsigned(9654, 14) & to_unsigned(6095, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    39 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(39, 6) & to_unsigned(14311, 14) & to_unsigned(7667, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    40 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(40, 6) & to_unsigned(15617, 14) & to_unsigned(8146, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    41 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(41, 6) & to_unsigned(4588, 14) & to_unsigned(11218, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    42 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(42, 6) & to_unsigned(13660, 14) & to_unsigned(6243, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    43 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(43, 6) & to_unsigned(8578, 14) & to_unsigned(7874, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    44 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(44, 6) & to_unsigned(11741, 14) & to_unsigned(2686, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    45 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(0, 6) & to_unsigned(1022, 14) & to_unsigned(1264, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    46 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1, 6) & to_unsigned(12604, 14) & to_unsigned(9965, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    47 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(2, 6) & to_unsigned(8217, 14) & to_unsigned(2707, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    48 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3, 6) & to_unsigned(3156, 14) & to_unsigned(11793, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    49 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 6) & to_unsigned(354, 14) & to_unsigned(1514, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    50 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 6) & to_unsigned(6978, 14) & to_unsigned(14058, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    51 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 6) & to_unsigned(7922, 14) & to_unsigned(16079, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    52 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 6) & to_unsigned(15087, 14) & to_unsigned(12138, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    53 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(8, 6) & to_unsigned(5053, 14) & to_unsigned(6470, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    54 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9, 6) & to_unsigned(12687, 14) & to_unsigned(14932, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    55 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10, 6) & to_unsigned(15458, 14) & to_unsigned(1763, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    56 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(11, 6) & to_unsigned(8121, 14) & to_unsigned(1721, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    57 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(12, 6) & to_unsigned(12431, 14) & to_unsigned(549, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    58 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(13, 6) & to_unsigned(4129, 14) & to_unsigned(7091, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    59 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(14, 6) & to_unsigned(1426, 14) & to_unsigned(8415, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    60 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(15, 6) & to_unsigned(9783, 14) & to_unsigned(7604, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    61 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(16, 6) & to_unsigned(6295, 14) & to_unsigned(11329, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    62 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(17, 6) & to_unsigned(1409, 14) & to_unsigned(12061, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    63 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(18, 6) & to_unsigned(8065, 14) & to_unsigned(9087, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    64 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(19, 6) & to_unsigned(2918, 14) & to_unsigned(8438, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    65 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(20, 6) & to_unsigned(1293, 14) & to_unsigned(14115, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    66 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(21, 6) & to_unsigned(3922, 14) & to_unsigned(13851, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    67 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(22, 6) & to_unsigned(3851, 14) & to_unsigned(4000, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    68 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(23, 6) & to_unsigned(5865, 14) & to_unsigned(1768, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    69 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(24, 6) & to_unsigned(2655, 14) & to_unsigned(14957, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    70 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(25, 6) & to_unsigned(5565, 14) & to_unsigned(6332, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    71 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(26, 6) & to_unsigned(4303, 14) & to_unsigned(12631, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    72 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(27, 6) & to_unsigned(11653, 14) & to_unsigned(12236, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    73 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(28, 6) & to_unsigned(16025, 14) & to_unsigned(7632, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    74 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(29, 6) & to_unsigned(4655, 14) & to_unsigned(14128, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    75 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(30, 6) & to_unsigned(9584, 14) & to_unsigned(13123, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    76 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(31, 6) & to_unsigned(13987, 14) & to_unsigned(9597, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    77 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(32, 6) & to_unsigned(15409, 14) & to_unsigned(12110, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    78 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(33, 6) & to_unsigned(8754, 14) & to_unsigned(15490, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    79 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(34, 6) & to_unsigned(7416, 14) & to_unsigned(15325, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    80 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(35, 6) & to_unsigned(2909, 14) & to_unsigned(15549, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    81 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(36, 6) & to_unsigned(2995, 14) & to_unsigned(8257, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    82 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(37, 6) & to_unsigned(9406, 14) & to_unsigned(4791, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    83 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(38, 6) & to_unsigned(11111, 14) & to_unsigned(4854, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    84 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(39, 6) & to_unsigned(2812, 14) & to_unsigned(8521, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    85 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(40, 6) & to_unsigned(8476, 14) & to_unsigned(14717, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    86 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(41, 6) & to_unsigned(7820, 14) & to_unsigned(15360, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    87 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(42, 6) & to_unsigned(1179, 14) & to_unsigned(7939, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    88 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(43, 6) & to_unsigned(2357, 14) & to_unsigned(8678, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    89 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(44, 6) & to_unsigned(7703, 14) & to_unsigned(6216, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    90 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(0, 6) & to_unsigned(3477, 14) & to_unsigned(7067, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    91 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1, 6) & to_unsigned(3931, 14) & to_unsigned(13845, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    92 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(2, 6) & to_unsigned(7675, 14) & to_unsigned(12899, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    93 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3, 6) & to_unsigned(1754, 14) & to_unsigned(8187, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    94 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 6) & to_unsigned(7785, 14) & to_unsigned(1400, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    95 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 6) & to_unsigned(9213, 14) & to_unsigned(5891, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    96 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 6) & to_unsigned(2494, 14) & to_unsigned(7703, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    97 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 6) & to_unsigned(2576, 14) & to_unsigned(7902, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    98 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(8, 6) & to_unsigned(4821, 14) & to_unsigned(15682, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    99 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9, 6) & to_unsigned(10426, 14) & to_unsigned(11935, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    100 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10, 6) & to_unsigned(1810, 14) & to_unsigned(904, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    101 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(11, 6) & to_unsigned(11332, 14) & to_unsigned(9264, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    102 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(12, 6) & to_unsigned(11312, 14) & to_unsigned(3570, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    103 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(13, 6) & to_unsigned(14916, 14) & to_unsigned(2650, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    104 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(14, 6) & to_unsigned(7679, 14) & to_unsigned(7842, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    105 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(15, 6) & to_unsigned(6089, 14) & to_unsigned(13084, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    106 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(16, 6) & to_unsigned(3938, 14) & to_unsigned(2751, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    107 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(17, 6) & to_unsigned(8509, 14) & to_unsigned(4648, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    108 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(18, 6) & to_unsigned(12204, 14) & to_unsigned(8917, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    109 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(19, 6) & to_unsigned(5749, 14) & to_unsigned(12443, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    110 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(20, 6) & to_unsigned(12613, 14) & to_unsigned(4431, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    111 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(21, 6) & to_unsigned(1344, 14) & to_unsigned(4014, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    112 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(22, 6) & to_unsigned(8488, 14) & to_unsigned(13850, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    113 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(23, 6) & to_unsigned(1730, 14) & to_unsigned(14896, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    114 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(24, 6) & to_unsigned(14942, 14) & to_unsigned(7126, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    115 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(25, 6) & to_unsigned(14983, 14) & to_unsigned(8863, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    116 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(26, 6) & to_unsigned(6578, 14) & to_unsigned(8564, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    117 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(27, 6) & to_unsigned(4947, 14) & to_unsigned(396, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    118 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(28, 6) & to_unsigned(297, 14) & to_unsigned(12805, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    119 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(29, 6) & to_unsigned(13878, 14) & to_unsigned(6692, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    120 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(30, 6) & to_unsigned(11857, 14) & to_unsigned(11186, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    121 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(31, 6) & to_unsigned(14395, 14) & to_unsigned(11493, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    122 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(32, 6) & to_unsigned(16145, 14) & to_unsigned(12251, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    123 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(33, 6) & to_unsigned(13462, 14) & to_unsigned(7428, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    124 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(34, 6) & to_unsigned(14526, 14) & to_unsigned(13119, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    125 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(35, 6) & to_unsigned(2535, 14) & to_unsigned(11243, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    126 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(36, 6) & to_unsigned(6465, 14) & to_unsigned(12690, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    127 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(37, 6) & to_unsigned(6872, 14) & to_unsigned(9334, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    128 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(38, 6) & to_unsigned(15371, 14) & to_unsigned(14023, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    129 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(39, 6) & to_unsigned(8101, 14) & to_unsigned(10187, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    130 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(40, 6) & to_unsigned(11963, 14) & to_unsigned(4848, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    131 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(41, 6) & to_unsigned(15125, 14) & to_unsigned(6119, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    132 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(42, 6) & to_unsigned(8051, 14) & to_unsigned(14465, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    133 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(43, 6) & to_unsigned(11139, 14) & to_unsigned(5167, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    134 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(44, 6) & to_unsigned(2883, 14) & to_unsigned(14521, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U'))
  );

  -- From /home/souto/phase4ground/tables/ldpc/dvb/orig/dvb_64800_s2_b8_t2_a5.txt, table is 144x150 (2700.0 bytes)
  -- Resource estimation: 9 x 18 kB BRAMs or 5 x 36 kB BRAMs
  type dvb_64800_s2_b8_t2_a5_t is array (143 downto 0) of std_logic_vector(149 downto 0);

  constant DVB_64800_S2_B8_T2_A5_COLUMN_WIDTHS : integer_array_t := (0 => 4, 1 => 6, 2 => 14, 3 => 14, 4 => 14, 5 => 14, 6 => 14, 7 => 14, 8 => 14, 9 => 14, 10 => 14, 11 => 14);

  constant DVB_64800_S2_B8_T2_A5 : dvb_64800_s2_b8_t2_a5_t := (
    0 => std_logic_vector(to_unsigned(11, 4) & to_unsigned(0, 6) & to_unsigned(149, 14) & to_unsigned(11212, 14) & to_unsigned(5575, 14) & to_unsigned(6360, 14) & to_unsigned(12559, 14) & to_unsigned(8108, 14) & to_unsigned(8505, 14) & to_unsigned(408, 14) & to_unsigned(10026, 14) & to_unsigned(12828, 14)),
    1 => std_logic_vector(to_unsigned(11, 4) & to_unsigned(1, 6) & to_unsigned(5237, 14) & to_unsigned(490, 14) & to_unsigned(10677, 14) & to_unsigned(4998, 14) & to_unsigned(3869, 14) & to_unsigned(3734, 14) & to_unsigned(3092, 14) & to_unsigned(3509, 14) & to_unsigned(7703, 14) & to_unsigned(10305, 14)),
    2 => std_logic_vector(to_unsigned(11, 4) & to_unsigned(2, 6) & to_unsigned(8742, 14) & to_unsigned(5553, 14) & to_unsigned(2820, 14) & to_unsigned(7085, 14) & to_unsigned(12116, 14) & to_unsigned(10485, 14) & to_unsigned(564, 14) & to_unsigned(7795, 14) & to_unsigned(2972, 14) & to_unsigned(2157, 14)),
    3 => std_logic_vector(to_unsigned(11, 4) & to_unsigned(3, 6) & to_unsigned(2699, 14) & to_unsigned(4304, 14) & to_unsigned(8350, 14) & to_unsigned(712, 14) & to_unsigned(2841, 14) & to_unsigned(3250, 14) & to_unsigned(4731, 14) & to_unsigned(10105, 14) & to_unsigned(517, 14) & to_unsigned(7516, 14)),
    4 => std_logic_vector(to_unsigned(11, 4) & to_unsigned(4, 6) & to_unsigned(12067, 14) & to_unsigned(1351, 14) & to_unsigned(11992, 14) & to_unsigned(12191, 14) & to_unsigned(11267, 14) & to_unsigned(5161, 14) & to_unsigned(537, 14) & to_unsigned(6166, 14) & to_unsigned(4246, 14) & to_unsigned(2363, 14)),
    5 => std_logic_vector(to_unsigned(11, 4) & to_unsigned(5, 6) & to_unsigned(6828, 14) & to_unsigned(7107, 14) & to_unsigned(2127, 14) & to_unsigned(3724, 14) & to_unsigned(5743, 14) & to_unsigned(11040, 14) & to_unsigned(10756, 14) & to_unsigned(4073, 14) & to_unsigned(1011, 14) & to_unsigned(3422, 14)),
    6 => std_logic_vector(to_unsigned(11, 4) & to_unsigned(6, 6) & to_unsigned(11259, 14) & to_unsigned(1216, 14) & to_unsigned(9526, 14) & to_unsigned(1466, 14) & to_unsigned(10816, 14) & to_unsigned(940, 14) & to_unsigned(3744, 14) & to_unsigned(2815, 14) & to_unsigned(11506, 14) & to_unsigned(11573, 14)),
    7 => std_logic_vector(to_unsigned(11, 4) & to_unsigned(7, 6) & to_unsigned(4549, 14) & to_unsigned(11507, 14) & to_unsigned(1118, 14) & to_unsigned(1274, 14) & to_unsigned(11751, 14) & to_unsigned(5207, 14) & to_unsigned(7854, 14) & to_unsigned(12803, 14) & to_unsigned(4047, 14) & to_unsigned(6484, 14)),
    8 => std_logic_vector(to_unsigned(11, 4) & to_unsigned(8, 6) & to_unsigned(8430, 14) & to_unsigned(4115, 14) & to_unsigned(9440, 14) & to_unsigned(413, 14) & to_unsigned(4455, 14) & to_unsigned(2262, 14) & to_unsigned(7915, 14) & to_unsigned(12402, 14) & to_unsigned(8579, 14) & to_unsigned(7052, 14)),
    9 => std_logic_vector(to_unsigned(11, 4) & to_unsigned(9, 6) & to_unsigned(3885, 14) & to_unsigned(9126, 14) & to_unsigned(5665, 14) & to_unsigned(4505, 14) & to_unsigned(2343, 14) & to_unsigned(253, 14) & to_unsigned(4707, 14) & to_unsigned(3742, 14) & to_unsigned(4166, 14) & to_unsigned(1556, 14)),
    10 => std_logic_vector(to_unsigned(11, 4) & to_unsigned(10, 6) & to_unsigned(1704, 14) & to_unsigned(8936, 14) & to_unsigned(6775, 14) & to_unsigned(8639, 14) & to_unsigned(8179, 14) & to_unsigned(7954, 14) & to_unsigned(8234, 14) & to_unsigned(7850, 14) & to_unsigned(8883, 14) & to_unsigned(8713, 14)),
    11 => std_logic_vector(to_unsigned(11, 4) & to_unsigned(11, 6) & to_unsigned(11716, 14) & to_unsigned(4344, 14) & to_unsigned(9087, 14) & to_unsigned(11264, 14) & to_unsigned(2274, 14) & to_unsigned(8832, 14) & to_unsigned(9147, 14) & to_unsigned(11930, 14) & to_unsigned(6054, 14) & to_unsigned(5455, 14)),
    12 => std_logic_vector(to_unsigned(11, 4) & to_unsigned(12, 6) & to_unsigned(7323, 14) & to_unsigned(3970, 14) & to_unsigned(10329, 14) & to_unsigned(2170, 14) & to_unsigned(8262, 14) & to_unsigned(3854, 14) & to_unsigned(2087, 14) & to_unsigned(12899, 14) & to_unsigned(9497, 14) & to_unsigned(11700, 14)),
    13 => std_logic_vector(to_unsigned(11, 4) & to_unsigned(13, 6) & to_unsigned(4418, 14) & to_unsigned(1467, 14) & to_unsigned(2490, 14) & to_unsigned(5841, 14) & to_unsigned(817, 14) & to_unsigned(11453, 14) & to_unsigned(533, 14) & to_unsigned(11217, 14) & to_unsigned(11962, 14) & to_unsigned(5251, 14)),
    14 => std_logic_vector(to_unsigned(11, 4) & to_unsigned(14, 6) & to_unsigned(1541, 14) & to_unsigned(4525, 14) & to_unsigned(7976, 14) & to_unsigned(3457, 14) & to_unsigned(9536, 14) & to_unsigned(7725, 14) & to_unsigned(3788, 14) & to_unsigned(2982, 14) & to_unsigned(6307, 14) & to_unsigned(5997, 14)),
    15 => std_logic_vector(to_unsigned(11, 4) & to_unsigned(15, 6) & to_unsigned(11484, 14) & to_unsigned(2739, 14) & to_unsigned(4023, 14) & to_unsigned(12107, 14) & to_unsigned(6516, 14) & to_unsigned(551, 14) & to_unsigned(2572, 14) & to_unsigned(6628, 14) & to_unsigned(8150, 14) & to_unsigned(9852, 14)),
    16 => std_logic_vector(to_unsigned(11, 4) & to_unsigned(16, 6) & to_unsigned(6070, 14) & to_unsigned(1761, 14) & to_unsigned(4627, 14) & to_unsigned(6534, 14) & to_unsigned(7913, 14) & to_unsigned(3730, 14) & to_unsigned(11866, 14) & to_unsigned(1813, 14) & to_unsigned(12306, 14) & to_unsigned(8249, 14)),
    17 => std_logic_vector(to_unsigned(11, 4) & to_unsigned(17, 6) & to_unsigned(12441, 14) & to_unsigned(5489, 14) & to_unsigned(8748, 14) & to_unsigned(7837, 14) & to_unsigned(7660, 14) & to_unsigned(2102, 14) & to_unsigned(11341, 14) & to_unsigned(2936, 14) & to_unsigned(6712, 14) & to_unsigned(11977, 14)),
    18 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(18, 6) & to_unsigned(10155, 14) & to_unsigned(4210, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    19 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(19, 6) & to_unsigned(1010, 14) & to_unsigned(10483, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    20 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(20, 6) & to_unsigned(8900, 14) & to_unsigned(10250, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    21 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(21, 6) & to_unsigned(10243, 14) & to_unsigned(12278, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    22 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(22, 6) & to_unsigned(7070, 14) & to_unsigned(4397, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    23 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(23, 6) & to_unsigned(12271, 14) & to_unsigned(3887, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    24 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(24, 6) & to_unsigned(11980, 14) & to_unsigned(6836, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    25 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(25, 6) & to_unsigned(9514, 14) & to_unsigned(4356, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    26 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(26, 6) & to_unsigned(7137, 14) & to_unsigned(10281, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    27 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(27, 6) & to_unsigned(11881, 14) & to_unsigned(2526, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    28 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(28, 6) & to_unsigned(1969, 14) & to_unsigned(11477, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    29 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(29, 6) & to_unsigned(3044, 14) & to_unsigned(10921, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    30 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(30, 6) & to_unsigned(2236, 14) & to_unsigned(8724, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    31 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(31, 6) & to_unsigned(9104, 14) & to_unsigned(6340, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    32 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(32, 6) & to_unsigned(7342, 14) & to_unsigned(8582, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    33 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(33, 6) & to_unsigned(11675, 14) & to_unsigned(10405, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    34 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(34, 6) & to_unsigned(6467, 14) & to_unsigned(12775, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    35 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(35, 6) & to_unsigned(3186, 14) & to_unsigned(12198, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    36 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(0, 6) & to_unsigned(9621, 14) & to_unsigned(11445, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    37 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1, 6) & to_unsigned(7486, 14) & to_unsigned(5611, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    38 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(2, 6) & to_unsigned(4319, 14) & to_unsigned(4879, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    39 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3, 6) & to_unsigned(2196, 14) & to_unsigned(344, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    40 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 6) & to_unsigned(7527, 14) & to_unsigned(6650, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    41 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 6) & to_unsigned(10693, 14) & to_unsigned(2440, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    42 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 6) & to_unsigned(6755, 14) & to_unsigned(2706, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    43 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 6) & to_unsigned(5144, 14) & to_unsigned(5998, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    44 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(8, 6) & to_unsigned(11043, 14) & to_unsigned(8033, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    45 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9, 6) & to_unsigned(4846, 14) & to_unsigned(4435, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    46 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10, 6) & to_unsigned(4157, 14) & to_unsigned(9228, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    47 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(11, 6) & to_unsigned(12270, 14) & to_unsigned(6562, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    48 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(12, 6) & to_unsigned(11954, 14) & to_unsigned(7592, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    49 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(13, 6) & to_unsigned(7420, 14) & to_unsigned(2592, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    50 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(14, 6) & to_unsigned(8810, 14) & to_unsigned(9636, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    51 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(15, 6) & to_unsigned(689, 14) & to_unsigned(5430, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    52 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(16, 6) & to_unsigned(920, 14) & to_unsigned(1304, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    53 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(17, 6) & to_unsigned(1253, 14) & to_unsigned(11934, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    54 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(18, 6) & to_unsigned(9559, 14) & to_unsigned(6016, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    55 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(19, 6) & to_unsigned(312, 14) & to_unsigned(7589, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    56 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(20, 6) & to_unsigned(4439, 14) & to_unsigned(4197, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    57 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(21, 6) & to_unsigned(4002, 14) & to_unsigned(9555, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    58 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(22, 6) & to_unsigned(12232, 14) & to_unsigned(7779, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    59 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(23, 6) & to_unsigned(1494, 14) & to_unsigned(8782, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    60 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(24, 6) & to_unsigned(10749, 14) & to_unsigned(3969, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    61 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(25, 6) & to_unsigned(4368, 14) & to_unsigned(3479, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    62 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(26, 6) & to_unsigned(6316, 14) & to_unsigned(5342, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    63 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(27, 6) & to_unsigned(2455, 14) & to_unsigned(3493, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    64 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(28, 6) & to_unsigned(12157, 14) & to_unsigned(7405, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    65 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(29, 6) & to_unsigned(6598, 14) & to_unsigned(11495, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    66 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(30, 6) & to_unsigned(11805, 14) & to_unsigned(4455, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    67 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(31, 6) & to_unsigned(9625, 14) & to_unsigned(2090, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    68 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(32, 6) & to_unsigned(4731, 14) & to_unsigned(2321, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    69 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(33, 6) & to_unsigned(3578, 14) & to_unsigned(2608, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    70 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(34, 6) & to_unsigned(8504, 14) & to_unsigned(1849, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    71 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(35, 6) & to_unsigned(4027, 14) & to_unsigned(1151, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    72 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(0, 6) & to_unsigned(5647, 14) & to_unsigned(4935, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    73 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1, 6) & to_unsigned(4219, 14) & to_unsigned(1870, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    74 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(2, 6) & to_unsigned(10968, 14) & to_unsigned(8054, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    75 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3, 6) & to_unsigned(6970, 14) & to_unsigned(5447, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    76 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 6) & to_unsigned(3217, 14) & to_unsigned(5638, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    77 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 6) & to_unsigned(8972, 14) & to_unsigned(669, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    78 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 6) & to_unsigned(5618, 14) & to_unsigned(12472, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    79 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 6) & to_unsigned(1457, 14) & to_unsigned(1280, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    80 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(8, 6) & to_unsigned(8868, 14) & to_unsigned(3883, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    81 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9, 6) & to_unsigned(8866, 14) & to_unsigned(1224, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    82 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10, 6) & to_unsigned(8371, 14) & to_unsigned(5972, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    83 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(11, 6) & to_unsigned(266, 14) & to_unsigned(4405, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    84 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(12, 6) & to_unsigned(3706, 14) & to_unsigned(3244, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    85 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(13, 6) & to_unsigned(6039, 14) & to_unsigned(5844, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    86 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(14, 6) & to_unsigned(7200, 14) & to_unsigned(3283, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    87 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(15, 6) & to_unsigned(1502, 14) & to_unsigned(11282, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    88 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(16, 6) & to_unsigned(12318, 14) & to_unsigned(2202, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    89 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(17, 6) & to_unsigned(4523, 14) & to_unsigned(965, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    90 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(18, 6) & to_unsigned(9587, 14) & to_unsigned(7011, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    91 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(19, 6) & to_unsigned(2552, 14) & to_unsigned(2051, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    92 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(20, 6) & to_unsigned(12045, 14) & to_unsigned(10306, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    93 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(21, 6) & to_unsigned(11070, 14) & to_unsigned(5104, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    94 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(22, 6) & to_unsigned(6627, 14) & to_unsigned(6906, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    95 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(23, 6) & to_unsigned(9889, 14) & to_unsigned(2121, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    96 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(24, 6) & to_unsigned(829, 14) & to_unsigned(9701, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    97 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(25, 6) & to_unsigned(2201, 14) & to_unsigned(1819, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    98 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(26, 6) & to_unsigned(6689, 14) & to_unsigned(12925, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    99 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(27, 6) & to_unsigned(2139, 14) & to_unsigned(8757, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    100 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(28, 6) & to_unsigned(12004, 14) & to_unsigned(5948, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    101 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(29, 6) & to_unsigned(8704, 14) & to_unsigned(3191, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    102 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(30, 6) & to_unsigned(8171, 14) & to_unsigned(10933, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    103 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(31, 6) & to_unsigned(6297, 14) & to_unsigned(7116, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    104 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(32, 6) & to_unsigned(616, 14) & to_unsigned(7146, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    105 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(33, 6) & to_unsigned(5142, 14) & to_unsigned(9761, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    106 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(34, 6) & to_unsigned(10377, 14) & to_unsigned(8138, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    107 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(35, 6) & to_unsigned(7616, 14) & to_unsigned(5811, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    108 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(0, 6) & to_unsigned(7285, 14) & to_unsigned(9863, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    109 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1, 6) & to_unsigned(7764, 14) & to_unsigned(10867, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    110 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(2, 6) & to_unsigned(12343, 14) & to_unsigned(9019, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    111 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3, 6) & to_unsigned(4414, 14) & to_unsigned(8331, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    112 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 6) & to_unsigned(3464, 14) & to_unsigned(642, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    113 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 6) & to_unsigned(6960, 14) & to_unsigned(2039, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    114 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 6) & to_unsigned(786, 14) & to_unsigned(3021, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    115 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 6) & to_unsigned(710, 14) & to_unsigned(2086, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    116 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(8, 6) & to_unsigned(7423, 14) & to_unsigned(5601, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    117 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9, 6) & to_unsigned(8120, 14) & to_unsigned(4885, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    118 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10, 6) & to_unsigned(12385, 14) & to_unsigned(11990, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    119 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(11, 6) & to_unsigned(9739, 14) & to_unsigned(10034, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    120 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(12, 6) & to_unsigned(424, 14) & to_unsigned(10162, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    121 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(13, 6) & to_unsigned(1347, 14) & to_unsigned(7597, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    122 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(14, 6) & to_unsigned(1450, 14) & to_unsigned(112, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    123 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(15, 6) & to_unsigned(7965, 14) & to_unsigned(8478, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    124 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(16, 6) & to_unsigned(8945, 14) & to_unsigned(7397, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    125 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(17, 6) & to_unsigned(6590, 14) & to_unsigned(8316, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    126 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(18, 6) & to_unsigned(6838, 14) & to_unsigned(9011, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    127 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(19, 6) & to_unsigned(6174, 14) & to_unsigned(9410, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    128 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(20, 6) & to_unsigned(255, 14) & to_unsigned(113, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    129 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(21, 6) & to_unsigned(6197, 14) & to_unsigned(5835, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    130 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(22, 6) & to_unsigned(12902, 14) & to_unsigned(3844, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    131 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(23, 6) & to_unsigned(4377, 14) & to_unsigned(3505, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    132 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(24, 6) & to_unsigned(5478, 14) & to_unsigned(8672, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    133 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(25, 6) & to_unsigned(4453, 14) & to_unsigned(2132, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    134 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(26, 6) & to_unsigned(9724, 14) & to_unsigned(1380, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    135 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(27, 6) & to_unsigned(12131, 14) & to_unsigned(11526, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    136 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(28, 6) & to_unsigned(12323, 14) & to_unsigned(9511, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    137 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(29, 6) & to_unsigned(8231, 14) & to_unsigned(1752, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    138 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(30, 6) & to_unsigned(497, 14) & to_unsigned(9022, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    139 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(31, 6) & to_unsigned(9288, 14) & to_unsigned(3080, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    140 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(32, 6) & to_unsigned(2481, 14) & to_unsigned(7515, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    141 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(33, 6) & to_unsigned(2696, 14) & to_unsigned(268, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    142 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(34, 6) & to_unsigned(4023, 14) & to_unsigned(12341, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    143 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(35, 6) & to_unsigned(7108, 14) & to_unsigned(5553, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U'))
  );

  -- From /home/souto/phase4ground/tables/ldpc/dvb/orig/dvb_64800_s2_b9_t2_a6.txt, table is 150x177 (3318.75 bytes)
  -- Resource estimation: 10 x 18 kB BRAMs or 5 x 36 kB BRAMs
  type dvb_64800_s2_b9_t2_a6_t is array (149 downto 0) of std_logic_vector(176 downto 0);

  constant DVB_64800_S2_B9_T2_A6_COLUMN_WIDTHS : integer_array_t := (0 => 4, 1 => 5, 2 => 14, 3 => 14, 4 => 14, 5 => 14, 6 => 14, 7 => 14, 8 => 14, 9 => 14, 10 => 14, 11 => 14, 12 => 14, 13 => 14);

  constant DVB_64800_S2_B9_T2_A6 : dvb_64800_s2_b9_t2_a6_t := (
    0 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(0, 5) & to_unsigned(4362, 14) & to_unsigned(416, 14) & to_unsigned(8909, 14) & to_unsigned(4156, 14) & to_unsigned(3216, 14) & to_unsigned(3112, 14) & to_unsigned(2560, 14) & to_unsigned(2912, 14) & to_unsigned(6405, 14) & to_unsigned(8593, 14) & to_unsigned(4969, 14) & to_unsigned(6723, 14)),
    1 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(1, 5) & to_unsigned(2479, 14) & to_unsigned(1786, 14) & to_unsigned(8978, 14) & to_unsigned(3011, 14) & to_unsigned(4339, 14) & to_unsigned(9313, 14) & to_unsigned(6397, 14) & to_unsigned(2957, 14) & to_unsigned(7288, 14) & to_unsigned(5484, 14) & to_unsigned(6031, 14) & to_unsigned(10217, 14)),
    2 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(2, 5) & to_unsigned(10175, 14) & to_unsigned(9009, 14) & to_unsigned(9889, 14) & to_unsigned(3091, 14) & to_unsigned(4985, 14) & to_unsigned(7267, 14) & to_unsigned(4092, 14) & to_unsigned(8874, 14) & to_unsigned(5671, 14) & to_unsigned(2777, 14) & to_unsigned(2189, 14) & to_unsigned(8716, 14)),
    3 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(3, 5) & to_unsigned(9052, 14) & to_unsigned(4795, 14) & to_unsigned(3924, 14) & to_unsigned(3370, 14) & to_unsigned(10058, 14) & to_unsigned(1128, 14) & to_unsigned(9996, 14) & to_unsigned(10165, 14) & to_unsigned(9360, 14) & to_unsigned(4297, 14) & to_unsigned(434, 14) & to_unsigned(5138, 14)),
    4 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(4, 5) & to_unsigned(2379, 14) & to_unsigned(7834, 14) & to_unsigned(4835, 14) & to_unsigned(2327, 14) & to_unsigned(9843, 14) & to_unsigned(804, 14) & to_unsigned(329, 14) & to_unsigned(8353, 14) & to_unsigned(7167, 14) & to_unsigned(3070, 14) & to_unsigned(1528, 14) & to_unsigned(7311, 14)),
    5 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(5, 5) & to_unsigned(3435, 14) & to_unsigned(7871, 14) & to_unsigned(348, 14) & to_unsigned(3693, 14) & to_unsigned(1876, 14) & to_unsigned(6585, 14) & to_unsigned(10340, 14) & to_unsigned(7144, 14) & to_unsigned(5870, 14) & to_unsigned(2084, 14) & to_unsigned(4052, 14) & to_unsigned(2780, 14)),
    6 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(6, 5) & to_unsigned(3917, 14) & to_unsigned(3111, 14) & to_unsigned(3476, 14) & to_unsigned(1304, 14) & to_unsigned(10331, 14) & to_unsigned(5939, 14) & to_unsigned(5199, 14) & to_unsigned(1611, 14) & to_unsigned(1991, 14) & to_unsigned(699, 14) & to_unsigned(8316, 14) & to_unsigned(9960, 14)),
    7 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(7, 5) & to_unsigned(6883, 14) & to_unsigned(3237, 14) & to_unsigned(1717, 14) & to_unsigned(10752, 14) & to_unsigned(7891, 14) & to_unsigned(9764, 14) & to_unsigned(4745, 14) & to_unsigned(3888, 14) & to_unsigned(10009, 14) & to_unsigned(4176, 14) & to_unsigned(4614, 14) & to_unsigned(1567, 14)),
    8 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(8, 5) & to_unsigned(10587, 14) & to_unsigned(2195, 14) & to_unsigned(1689, 14) & to_unsigned(2968, 14) & to_unsigned(5420, 14) & to_unsigned(2580, 14) & to_unsigned(2883, 14) & to_unsigned(6496, 14) & to_unsigned(111, 14) & to_unsigned(6023, 14) & to_unsigned(1024, 14) & to_unsigned(4449, 14)),
    9 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(9, 5) & to_unsigned(3786, 14) & to_unsigned(8593, 14) & to_unsigned(2074, 14) & to_unsigned(3321, 14) & to_unsigned(5057, 14) & to_unsigned(1450, 14) & to_unsigned(3840, 14) & to_unsigned(5444, 14) & to_unsigned(6572, 14) & to_unsigned(3094, 14) & to_unsigned(9892, 14) & to_unsigned(1512, 14)),
    10 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(10, 5) & to_unsigned(8548, 14) & to_unsigned(1848, 14) & to_unsigned(10372, 14) & to_unsigned(4585, 14) & to_unsigned(7313, 14) & to_unsigned(6536, 14) & to_unsigned(6379, 14) & to_unsigned(1766, 14) & to_unsigned(9462, 14) & to_unsigned(2456, 14) & to_unsigned(5606, 14) & to_unsigned(9975, 14)),
    11 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(11, 5) & to_unsigned(8204, 14) & to_unsigned(10593, 14) & to_unsigned(7935, 14) & to_unsigned(3636, 14) & to_unsigned(3882, 14) & to_unsigned(394, 14) & to_unsigned(5968, 14) & to_unsigned(8561, 14) & to_unsigned(2395, 14) & to_unsigned(7289, 14) & to_unsigned(9267, 14) & to_unsigned(9978, 14)),
    12 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(12, 5) & to_unsigned(7795, 14) & to_unsigned(74, 14) & to_unsigned(1633, 14) & to_unsigned(9542, 14) & to_unsigned(6867, 14) & to_unsigned(7352, 14) & to_unsigned(6417, 14) & to_unsigned(7568, 14) & to_unsigned(10623, 14) & to_unsigned(725, 14) & to_unsigned(2531, 14) & to_unsigned(9115, 14)),
    13 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(13, 5) & to_unsigned(7151, 14) & to_unsigned(2482, 14) & to_unsigned(4260, 14) & to_unsigned(5003, 14) & to_unsigned(10105, 14) & to_unsigned(7419, 14) & to_unsigned(9203, 14) & to_unsigned(6691, 14) & to_unsigned(8798, 14) & to_unsigned(2092, 14) & to_unsigned(8263, 14) & to_unsigned(3755, 14)),
    14 => std_logic_vector(to_unsigned(13, 4) & to_unsigned(14, 5) & to_unsigned(3600, 14) & to_unsigned(570, 14) & to_unsigned(4527, 14) & to_unsigned(200, 14) & to_unsigned(9718, 14) & to_unsigned(6771, 14) & to_unsigned(1995, 14) & to_unsigned(8902, 14) & to_unsigned(5446, 14) & to_unsigned(768, 14) & to_unsigned(1103, 14) & to_unsigned(6520, 14)),
    15 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(15, 5) & to_unsigned(6304, 14) & to_unsigned(7621, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    16 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(16, 5) & to_unsigned(6498, 14) & to_unsigned(9209, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    17 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(17, 5) & to_unsigned(7293, 14) & to_unsigned(6786, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    18 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(18, 5) & to_unsigned(5950, 14) & to_unsigned(1708, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    19 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(19, 5) & to_unsigned(8521, 14) & to_unsigned(1793, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    20 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(20, 5) & to_unsigned(6174, 14) & to_unsigned(7854, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    21 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(21, 5) & to_unsigned(9773, 14) & to_unsigned(1190, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    22 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(22, 5) & to_unsigned(9517, 14) & to_unsigned(10268, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    23 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(23, 5) & to_unsigned(2181, 14) & to_unsigned(9349, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    24 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(24, 5) & to_unsigned(1949, 14) & to_unsigned(5560, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    25 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(25, 5) & to_unsigned(1556, 14) & to_unsigned(555, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    26 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(26, 5) & to_unsigned(8600, 14) & to_unsigned(3827, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    27 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(27, 5) & to_unsigned(5072, 14) & to_unsigned(1057, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    28 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(28, 5) & to_unsigned(7928, 14) & to_unsigned(3542, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    29 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(29, 5) & to_unsigned(3226, 14) & to_unsigned(3762, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    30 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(0, 5) & to_unsigned(7045, 14) & to_unsigned(2420, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    31 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1, 5) & to_unsigned(9645, 14) & to_unsigned(2641, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    32 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(2, 5) & to_unsigned(2774, 14) & to_unsigned(2452, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    33 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3, 5) & to_unsigned(5331, 14) & to_unsigned(2031, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    34 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 5) & to_unsigned(9400, 14) & to_unsigned(7503, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    35 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 5) & to_unsigned(1850, 14) & to_unsigned(2338, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    36 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 5) & to_unsigned(10456, 14) & to_unsigned(9774, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    37 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 5) & to_unsigned(1692, 14) & to_unsigned(9276, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    38 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(8, 5) & to_unsigned(10037, 14) & to_unsigned(4038, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    39 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9, 5) & to_unsigned(3964, 14) & to_unsigned(338, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    40 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10, 5) & to_unsigned(2640, 14) & to_unsigned(5087, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    41 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(11, 5) & to_unsigned(858, 14) & to_unsigned(3473, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    42 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(12, 5) & to_unsigned(5582, 14) & to_unsigned(5683, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    43 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(13, 5) & to_unsigned(9523, 14) & to_unsigned(916, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    44 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(14, 5) & to_unsigned(4107, 14) & to_unsigned(1559, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    45 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(15, 5) & to_unsigned(4506, 14) & to_unsigned(3491, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    46 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(16, 5) & to_unsigned(8191, 14) & to_unsigned(4182, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    47 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(17, 5) & to_unsigned(10192, 14) & to_unsigned(6157, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    48 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(18, 5) & to_unsigned(5668, 14) & to_unsigned(3305, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    49 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(19, 5) & to_unsigned(3449, 14) & to_unsigned(1540, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    50 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(20, 5) & to_unsigned(4766, 14) & to_unsigned(2697, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    51 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(21, 5) & to_unsigned(4069, 14) & to_unsigned(6675, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    52 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(22, 5) & to_unsigned(1117, 14) & to_unsigned(1016, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    53 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(23, 5) & to_unsigned(5619, 14) & to_unsigned(3085, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    54 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(24, 5) & to_unsigned(8483, 14) & to_unsigned(8400, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    55 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(25, 5) & to_unsigned(8255, 14) & to_unsigned(394, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    56 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(26, 5) & to_unsigned(6338, 14) & to_unsigned(5042, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    57 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(27, 5) & to_unsigned(6174, 14) & to_unsigned(5119, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    58 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(28, 5) & to_unsigned(7203, 14) & to_unsigned(1989, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    59 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(29, 5) & to_unsigned(1781, 14) & to_unsigned(5174, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    60 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(0, 5) & to_unsigned(1464, 14) & to_unsigned(3559, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    61 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1, 5) & to_unsigned(3376, 14) & to_unsigned(4214, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    62 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(2, 5) & to_unsigned(7238, 14) & to_unsigned(67, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    63 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3, 5) & to_unsigned(10595, 14) & to_unsigned(8831, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    64 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 5) & to_unsigned(1221, 14) & to_unsigned(6513, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    65 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 5) & to_unsigned(5300, 14) & to_unsigned(4652, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    66 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 5) & to_unsigned(1429, 14) & to_unsigned(9749, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    67 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 5) & to_unsigned(7878, 14) & to_unsigned(5131, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    68 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(8, 5) & to_unsigned(4435, 14) & to_unsigned(10284, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    69 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9, 5) & to_unsigned(6331, 14) & to_unsigned(5507, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    70 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10, 5) & to_unsigned(6662, 14) & to_unsigned(4941, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    71 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(11, 5) & to_unsigned(9614, 14) & to_unsigned(10238, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    72 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(12, 5) & to_unsigned(8400, 14) & to_unsigned(8025, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    73 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(13, 5) & to_unsigned(9156, 14) & to_unsigned(5630, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    74 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(14, 5) & to_unsigned(7067, 14) & to_unsigned(8878, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    75 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(15, 5) & to_unsigned(9027, 14) & to_unsigned(3415, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    76 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(16, 5) & to_unsigned(1690, 14) & to_unsigned(3866, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    77 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(17, 5) & to_unsigned(2854, 14) & to_unsigned(8469, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    78 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(18, 5) & to_unsigned(6206, 14) & to_unsigned(630, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    79 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(19, 5) & to_unsigned(363, 14) & to_unsigned(5453, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    80 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(20, 5) & to_unsigned(4125, 14) & to_unsigned(7008, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    81 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(21, 5) & to_unsigned(1612, 14) & to_unsigned(6702, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    82 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(22, 5) & to_unsigned(9069, 14) & to_unsigned(9226, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    83 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(23, 5) & to_unsigned(5767, 14) & to_unsigned(4060, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    84 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(24, 5) & to_unsigned(3743, 14) & to_unsigned(9237, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    85 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(25, 5) & to_unsigned(7018, 14) & to_unsigned(5572, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    86 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(26, 5) & to_unsigned(8892, 14) & to_unsigned(4536, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    87 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(27, 5) & to_unsigned(853, 14) & to_unsigned(6064, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    88 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(28, 5) & to_unsigned(8069, 14) & to_unsigned(5893, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    89 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(29, 5) & to_unsigned(2051, 14) & to_unsigned(2885, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    90 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(0, 5) & to_unsigned(10691, 14) & to_unsigned(3153, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    91 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1, 5) & to_unsigned(3602, 14) & to_unsigned(4055, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    92 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(2, 5) & to_unsigned(328, 14) & to_unsigned(1717, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    93 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3, 5) & to_unsigned(2219, 14) & to_unsigned(9299, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    94 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 5) & to_unsigned(1939, 14) & to_unsigned(7898, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    95 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 5) & to_unsigned(617, 14) & to_unsigned(206, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    96 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 5) & to_unsigned(8544, 14) & to_unsigned(1374, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    97 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 5) & to_unsigned(10676, 14) & to_unsigned(3240, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    98 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(8, 5) & to_unsigned(6672, 14) & to_unsigned(9489, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    99 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9, 5) & to_unsigned(3170, 14) & to_unsigned(7457, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    100 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10, 5) & to_unsigned(7868, 14) & to_unsigned(5731, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    101 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(11, 5) & to_unsigned(6121, 14) & to_unsigned(10732, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    102 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(12, 5) & to_unsigned(4843, 14) & to_unsigned(9132, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    103 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(13, 5) & to_unsigned(580, 14) & to_unsigned(9591, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    104 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(14, 5) & to_unsigned(6267, 14) & to_unsigned(9290, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    105 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(15, 5) & to_unsigned(3009, 14) & to_unsigned(2268, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    106 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(16, 5) & to_unsigned(195, 14) & to_unsigned(2419, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    107 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(17, 5) & to_unsigned(8016, 14) & to_unsigned(1557, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    108 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(18, 5) & to_unsigned(1516, 14) & to_unsigned(9195, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    109 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(19, 5) & to_unsigned(8062, 14) & to_unsigned(9064, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    110 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(20, 5) & to_unsigned(2095, 14) & to_unsigned(8968, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    111 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(21, 5) & to_unsigned(753, 14) & to_unsigned(7326, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    112 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(22, 5) & to_unsigned(6291, 14) & to_unsigned(3833, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    113 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(23, 5) & to_unsigned(2614, 14) & to_unsigned(7844, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    114 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(24, 5) & to_unsigned(2303, 14) & to_unsigned(646, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    115 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(25, 5) & to_unsigned(2075, 14) & to_unsigned(611, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    116 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(26, 5) & to_unsigned(4687, 14) & to_unsigned(362, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    117 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(27, 5) & to_unsigned(8684, 14) & to_unsigned(9940, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    118 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(28, 5) & to_unsigned(4830, 14) & to_unsigned(2065, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    119 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(29, 5) & to_unsigned(7038, 14) & to_unsigned(1363, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    120 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(0, 5) & to_unsigned(1769, 14) & to_unsigned(7837, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    121 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(1, 5) & to_unsigned(3801, 14) & to_unsigned(1689, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    122 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(2, 5) & to_unsigned(10070, 14) & to_unsigned(2359, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    123 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(3, 5) & to_unsigned(3667, 14) & to_unsigned(9918, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    124 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(4, 5) & to_unsigned(1914, 14) & to_unsigned(6920, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    125 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(5, 5) & to_unsigned(4244, 14) & to_unsigned(5669, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    126 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(6, 5) & to_unsigned(10245, 14) & to_unsigned(7821, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    127 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(7, 5) & to_unsigned(7648, 14) & to_unsigned(3944, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    128 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(8, 5) & to_unsigned(3310, 14) & to_unsigned(5488, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    129 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(9, 5) & to_unsigned(6346, 14) & to_unsigned(9666, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    130 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(10, 5) & to_unsigned(7088, 14) & to_unsigned(6122, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    131 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(11, 5) & to_unsigned(1291, 14) & to_unsigned(7827, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    132 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(12, 5) & to_unsigned(10592, 14) & to_unsigned(8945, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    133 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(13, 5) & to_unsigned(3609, 14) & to_unsigned(7120, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    134 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(14, 5) & to_unsigned(9168, 14) & to_unsigned(9112, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    135 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(15, 5) & to_unsigned(6203, 14) & to_unsigned(8052, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    136 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(16, 5) & to_unsigned(3330, 14) & to_unsigned(2895, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    137 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(17, 5) & to_unsigned(4264, 14) & to_unsigned(10563, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    138 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(18, 5) & to_unsigned(10556, 14) & to_unsigned(6496, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    139 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(19, 5) & to_unsigned(8807, 14) & to_unsigned(7645, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    140 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(20, 5) & to_unsigned(1999, 14) & to_unsigned(4530, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    141 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(21, 5) & to_unsigned(9202, 14) & to_unsigned(6818, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    142 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(22, 5) & to_unsigned(3403, 14) & to_unsigned(1734, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    143 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(23, 5) & to_unsigned(2106, 14) & to_unsigned(9023, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    144 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(24, 5) & to_unsigned(6881, 14) & to_unsigned(3883, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    145 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(25, 5) & to_unsigned(3895, 14) & to_unsigned(2171, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    146 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(26, 5) & to_unsigned(4062, 14) & to_unsigned(6424, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    147 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(27, 5) & to_unsigned(3755, 14) & to_unsigned(9536, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    148 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(28, 5) & to_unsigned(4683, 14) & to_unsigned(2131, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U')),
    149 => std_logic_vector(to_unsigned(3, 4) & to_unsigned(29, 5) & to_unsigned(7347, 14) & to_unsigned(8027, 14) & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U') & (13 downto 0 => 'U'))
  );


end package ldpc_tables_pkg;

package body ldpc_tables_pkg is
end package body ldpc_tables_pkg;